module gameover(G,A,M,E,O,V,E2,R,clk,pixel_row,pixel_col);

input clk;
input [10:0]pixel_row,pixel_col;
output reg G,A,M,E,O,V,E2,R;

reg [39:0] line_G01,line_G02,line_G03,line_G04,line_G05,line_G06,line_G07,line_G08,line_G09,line_G10,line_G11,line_G12,line_G13,line_G14,line_G15;
reg [39:0] line_A01,line_A02,line_A03,line_A04,line_A05,line_A06,line_A07,line_A08,line_A09,line_A10,line_A11,line_A12,line_A13,line_A14,line_A15;
reg [39:0] line_M01,line_M02,line_M03,line_M04,line_M05,line_M06,line_M07,line_M08,line_M09,line_M10,line_M11,line_M12,line_M13,line_M14,line_M15;
reg [39:0] line_E01,line_E02,line_E03,line_E04,line_E05,line_E06,line_E07,line_E08,line_E09,line_E10,line_E11,line_E12,line_E13,line_E14,line_E15;
reg [39:0] line_O01,line_O02,line_O03,line_O04,line_O05,line_O06,line_O07,line_O08,line_O09,line_O10,line_O11,line_O12,line_O13,line_O14,line_O15;
reg [39:0] line_V01,line_V02,line_V03,line_V04,line_V05,line_V06,line_V07,line_V08,line_V09,line_V10,line_V11,line_V12,line_V13,line_V14,line_V15;
reg [39:0] line_R01,line_R02,line_R03,line_R04,line_R05,line_R06,line_R07,line_R08,line_R09,line_R10,line_R11,line_R12,line_R13,line_R14,line_R15;


always @(posedge clk) begin
		line_G01 <= 40'b0000000000000000000000000000000000000000;
		line_G02 <= 40'b0000000000000011111111111111111100000000;
		line_G03 <= 40'b0000000001111111111111111111111111100000;
		line_G04 <= 40'b0000000111111111000000000000000111100000;
		line_G05 <= 40'b0000011111111100000000000000000000000000;
		line_G06 <= 40'b0000111111110000000000000000000000000000;
		line_G07 <= 40'b0000111111100000000011111111111111000000;
		line_G08 <= 40'b0000111111100000000111111111111111100000;
		line_G09 <= 40'b0000111111110000000000000001111111100000;
		line_G09 <= 40'b0000011111111000000000000001111111100000;
		line_G10 <= 40'b0000001111111110000000000001111111100000;
		line_G11 <= 40'b0000000011111111111111111111111111100000;
		line_G12 <= 40'b0000000000111111111111111111111111000000;
		line_G14 <= 40'b0000000000000000001111111000000000000000;
		line_G15 <= 40'b0000000000000000000000000000000000000000;
end

always @(posedge clk) begin
		line_A01 <= 40'b0000000000000000000000000000000000000000;
		line_A02 <= 40'b0000000000000000111111111000000000000000;
		line_A03 <= 40'b0000000000000011111111111100000000000000;
		line_A04 <= 40'b0000000000000111111111111110000000000000;
		line_A05 <= 40'b0000000000001111111001111111000000000000;
		line_A06 <= 40'b0000000000011111110000111111100000000000;
		line_A07 <= 40'b0000000000111111100000011111110000000000;
		line_A08 <= 40'b0000000001111111000000001111111000000000;
		line_A09 <= 40'b0000000011111110000000000111111100000000;
		line_A09 <= 40'b0000000011111111111111111111111110000000;
		line_A10 <= 40'b0000001111111111111111111111111111000000;
		line_A11 <= 40'b0000011111110000000000000000111111100000;
		line_A12 <= 40'b0000111111100000000000000000011111110000;
		line_A14 <= 40'b0000111111000000000000000000001111111000;
		line_A15 <= 40'b0000000000000000000000000000000000000000;
end

always @(posedge clk) begin
		line_M01 <= 40'b0000000000000000000000000000000000000000;
		line_M02 <= 40'b0000000000000000000000000000000000000000;
		line_M03 <= 40'b1111111111110000000000000000011111111111;
		line_M04 <= 40'b1111111111111000000000000000111111111111;
		line_M05 <= 40'b1111110111111100000000000001111110011111;
		line_M06 <= 40'b1111110011111110000000000011111100011111;
		line_M07 <= 40'b1111110001111111000000000111111000011111;
		line_M08 <= 40'b1111110000111111100000001111110000011111;
		line_M09 <= 40'b1111110000011111110000011111100000011111;
		line_M09 <= 40'b1111110000001111111000111111000000011111;
		line_M10 <= 40'b1111110000000111111111111110000000011111;
		line_M11 <= 40'b1111110000000011111111111100000000011111;
		line_M12 <= 40'b1111110000000001111111111000000000011111;
		line_M14 <= 40'b1111110000000000111111110000000000011111;
		line_M15 <= 40'b0000000000000000000000000000000000000000;
end

always @(posedge clk) begin
		line_E01 <= 40'b0000000000000000000000000000000000000000;
		line_E02 <= 40'b0000000000000000000000000000000000000000;
		line_E03 <= 40'b0000000011111111111111111111100000000000;
		line_E04 <= 40'b0000000011111110000000000000000000000000;
		line_E05 <= 40'b0000000011111110000000000000000000000000;
		line_E06 <= 40'b0000000011111110000000000000000000000000;
		line_E07 <= 40'b0000000011111110000000000000000000000000;
		line_E08 <= 40'b0000000011111111111111111110000000000000;
		line_E09 <= 40'b0000000011111110000000000000000000000000;
		line_E09 <= 40'b0000000011111110000000000000000000000000;
		line_E10 <= 40'b0000000011111110000000000000000000000000;
		line_E11 <= 40'b0000000011111100000000000000000000000000;
		line_E12 <= 40'b0000000011111111111111111111100000000000;
		line_E14 <= 40'b0000000011111111111111111111100000000000;
		line_E15 <= 40'b0000000000000000000000000000000000000000;
end

always @(posedge clk) begin
		line_O01 <= 40'b0000000000000000000000000000000000000000;
		line_O02 <= 40'b0000000000000000011111111000000000000000;
		line_O03 <= 40'b0000000000111111111111111111111100000000;
		line_O04 <= 40'b0000000111111111100000001111111111100000;
		line_O05 <= 40'b0000011111111100000000000000111111110000;
		line_O06 <= 40'b0000111111110000000000000000011111111000;
		line_O07 <= 40'b0000111111100000000000000000001111111100;
		line_O08 <= 40'b0001111111100000000000000000001111111100;
		line_O09 <= 40'b0001111111100000000000000000001111111100;
		line_O09 <= 40'b0000111111110000000000000000001111111000;
		line_O10 <= 40'b0000111111111000000000000000111111110000;
		line_O11 <= 40'b0000001111111110000000000011111111100000;
		line_O12 <= 40'b0000000001111111111111111111111110000000;
		line_O14 <= 40'b0000000000001111111111111111000000000000;
		line_O15 <= 40'b0000000000000000000000000000000000000000;
end

always @(posedge clk) begin
		line_V01 <= 40'b0000000000000000000000000000000000000000;
		line_V02 <= 40'b0000111111100000000000000000001111110000;
		line_V03 <= 40'b0000111111110000000000000000011111110000;
		line_V04 <= 40'b0000001111111000000000000000111111100000;
		line_V05 <= 40'b0000000111111100000000000001111111000000;
		line_V06 <= 40'b0000000011111110000000000011111110000000;
		line_V07 <= 40'b0000000001111111000000000111111100000000;
		line_V08 <= 40'b0000000000111111100000001111111000000000;
		line_V09 <= 40'b0000000000011111110000011111110000000000;
		line_V09 <= 40'b0000000000001111111000111111100000000000;
		line_V10 <= 40'b0000000000000111111101111111000000000000;
		line_V11 <= 40'b0000000000000011111111111110000000000000;
		line_V12 <= 40'b0000000000000001111111111100000000000000;
		line_V14 <= 40'b0000000000000000111111110000000000000000;
		line_V15 <= 40'b0000000000000000000000000000000000000000;
end

always @(posedge clk) begin
		line_R01 <= 40'b0000000000000000000000000000000000000000;
		line_R02 <= 40'b0000000011111111111111110000000000000000;
		line_R03 <= 40'b0000000111111111111111111111100000000000;
		line_R04 <= 40'b0000000111111100000000111111111000000000;
		line_R05 <= 40'b0000000111111100000000001111111100000000;
		line_R06 <= 40'b0000000111111100000000001111111100000000;
		line_R07 <= 40'b0000000111111100000000111111111000000000;
		line_R08 <= 40'b0000000111111111111111111110000000000000;
		line_R09 <= 40'b0000000111111111111111111110000000000000;
		line_R09 <= 40'b0000000111111100000001111111100000000000;
		line_R10 <= 40'b0000000111111100000000011111110000000000;
		line_R11 <= 40'b0000000111111100000000001111111100000000;
		line_R12 <= 40'b0000000111111100000000000111111110000000;
		line_R14 <= 40'b0000000111111100000000000011111100000000;
		line_R15 <= 40'b0000000000000000000000000000000000000000;
end

always @(posedge clk) begin
	case (pixel_row)
		11'd323:
			case (pixel_col)
				11'd409:G <= line_G01[39];	11'd419:G <= line_G01[29];	11'd429:G <= line_G01[19];	11'd439:G <= line_G01[9];
				11'd410:G <= line_G01[38];	11'd420:G <= line_G01[28];	11'd430:G <= line_G01[18];	11'd440:G <= line_G01[8];
				11'd411:G <= line_G01[37];	11'd421:G <= line_G01[27];	11'd431:G <= line_G01[17];	11'd441:G <= line_G01[7];
				11'd412:G <= line_G01[36];	11'd422:G <= line_G01[26];	11'd432:G <= line_G01[16];	11'd442:G <= line_G01[6];
				11'd413:G <= line_G01[35];	11'd423:G <= line_G01[25];	11'd433:G <= line_G01[15];	11'd443:G <= line_G01[5];
				11'd414:G <= line_G01[34];	11'd424:G <= line_G01[24];	11'd434:G <= line_G01[14];	11'd444:G <= line_G01[4];
				11'd415:G <= line_G01[33];	11'd425:G <= line_G01[23];	11'd435:G <= line_G01[13];	11'd445:G <= line_G01[3];
				11'd416:G <= line_G01[32];	11'd426:G <= line_G01[22];	11'd436:G <= line_G01[12];	11'd446:G <= line_G01[2];
				11'd417:G <= line_G01[31];	11'd427:G <= line_G01[21];	11'd437:G <= line_G01[11];	11'd447:G <= line_G01[1];
				11'd418:G <= line_G01[30];	11'd428:G <= line_G01[20];	11'd438:G <= line_G01[10];	11'd448:G <= line_G01[0];
				default:G <= 0;
			endcase
		11'd324:
			case (pixel_col)
				11'd409:G <= line_G02[39];	11'd419:G <= line_G02[29];	11'd429:G <= line_G02[19];	11'd439:G <= line_G02[9];
				11'd410:G <= line_G02[38];	11'd420:G <= line_G02[28];	11'd430:G <= line_G02[18];	11'd440:G <= line_G02[8];
				11'd411:G <= line_G02[37];	11'd421:G <= line_G02[27];	11'd431:G <= line_G02[17];	11'd441:G <= line_G02[7];
				11'd412:G <= line_G02[36];	11'd422:G <= line_G02[26];	11'd432:G <= line_G02[16];	11'd442:G <= line_G02[6];
				11'd413:G <= line_G02[35];	11'd423:G <= line_G02[25];	11'd433:G <= line_G02[15];	11'd443:G <= line_G02[5];
				11'd414:G <= line_G02[34];	11'd424:G <= line_G02[24];	11'd434:G <= line_G02[14];	11'd444:G <= line_G02[4];
				11'd415:G <= line_G02[33];	11'd425:G <= line_G02[23];	11'd435:G <= line_G02[13];	11'd445:G <= line_G02[3];
				11'd416:G <= line_G02[32];	11'd426:G <= line_G02[22];	11'd436:G <= line_G02[12];	11'd446:G <= line_G02[2];
				11'd417:G <= line_G02[31];	11'd427:G <= line_G02[21];	11'd437:G <= line_G02[11];	11'd447:G <= line_G02[1];
				11'd418:G <= line_G02[30];	11'd428:G <= line_G02[20];	11'd438:G <= line_G02[10];	11'd448:G <= line_G02[0];
				default:G <= 0;
			endcase
		11'd325:
			case (pixel_col)
				11'd409:G <= line_G03[39];	11'd419:G <= line_G03[29];	11'd429:G <= line_G03[19];	11'd439:G <= line_G03[9];
				11'd410:G <= line_G03[38];	11'd420:G <= line_G03[28];	11'd430:G <= line_G03[18];	11'd440:G <= line_G03[8];
				11'd411:G <= line_G03[37];	11'd421:G <= line_G03[27];	11'd431:G <= line_G03[17];	11'd441:G <= line_G03[7];
				11'd412:G <= line_G03[36];	11'd422:G <= line_G03[26];	11'd432:G <= line_G03[16];	11'd442:G <= line_G03[6];
				11'd413:G <= line_G03[35];	11'd423:G <= line_G03[25];	11'd433:G <= line_G03[15];	11'd443:G <= line_G03[5];
				11'd414:G <= line_G03[34];	11'd424:G <= line_G03[24];	11'd434:G <= line_G03[14];	11'd444:G <= line_G03[4];
				11'd415:G <= line_G03[33];	11'd425:G <= line_G03[23];	11'd435:G <= line_G03[13];	11'd445:G <= line_G03[3];
				11'd416:G <= line_G03[32];	11'd426:G <= line_G03[22];	11'd436:G <= line_G03[12];	11'd446:G <= line_G03[2];
				11'd417:G <= line_G03[31];	11'd427:G <= line_G03[21];	11'd437:G <= line_G03[11];	11'd447:G <= line_G03[1];
				11'd418:G <= line_G03[30];	11'd428:G <= line_G03[20];	11'd438:G <= line_G03[10];	11'd448:G <= line_G03[0];
				default:G <= 0;
			endcase
		11'd326:
			case (pixel_col)
				11'd409:G <= line_G04[39];	11'd419:G <= line_G04[29];	11'd429:G <= line_G04[19];	11'd439:G <= line_G04[9];
				11'd410:G <= line_G04[38];	11'd420:G <= line_G04[28];	11'd430:G <= line_G04[18];	11'd440:G <= line_G04[8];
				11'd411:G <= line_G04[37];	11'd421:G <= line_G04[27];	11'd431:G <= line_G04[17];	11'd441:G <= line_G04[7];
				11'd412:G <= line_G04[36];	11'd422:G <= line_G04[26];	11'd432:G <= line_G04[16];	11'd442:G <= line_G04[6];
				11'd413:G <= line_G04[35];	11'd423:G <= line_G04[25];	11'd433:G <= line_G04[15];	11'd443:G <= line_G04[5];
				11'd414:G <= line_G04[34];	11'd424:G <= line_G04[24];	11'd434:G <= line_G04[14];	11'd444:G <= line_G04[4];
				11'd415:G <= line_G04[33];	11'd425:G <= line_G04[23];	11'd435:G <= line_G04[13];	11'd445:G <= line_G04[3];
				11'd416:G <= line_G04[32];	11'd426:G <= line_G04[22];	11'd436:G <= line_G04[12];	11'd446:G <= line_G04[2];
				11'd417:G <= line_G04[31];	11'd427:G <= line_G04[21];	11'd437:G <= line_G04[11];	11'd447:G <= line_G04[1];
				11'd418:G <= line_G04[30];	11'd428:G <= line_G04[20];	11'd438:G <= line_G04[10];	11'd448:G <= line_G04[0];
				default:G <= 0;
			endcase
		11'd327:
			case (pixel_col)
				11'd409:G <= line_G05[39];	11'd419:G <= line_G05[29];	11'd429:G <= line_G05[19];	11'd439:G <= line_G05[9];
				11'd410:G <= line_G05[38];	11'd420:G <= line_G05[28];	11'd430:G <= line_G05[18];	11'd440:G <= line_G05[8];
				11'd411:G <= line_G05[37];	11'd421:G <= line_G05[27];	11'd431:G <= line_G05[17];	11'd441:G <= line_G05[7];
				11'd412:G <= line_G05[36];	11'd422:G <= line_G05[26];	11'd432:G <= line_G05[16];	11'd442:G <= line_G05[6];
				11'd413:G <= line_G05[35];	11'd423:G <= line_G05[25];	11'd433:G <= line_G05[15];	11'd443:G <= line_G05[5];
				11'd414:G <= line_G05[34];	11'd424:G <= line_G05[24];	11'd434:G <= line_G05[14];	11'd444:G <= line_G05[4];
				11'd415:G <= line_G05[33];	11'd425:G <= line_G05[23];	11'd435:G <= line_G05[13];	11'd445:G <= line_G05[3];
				11'd416:G <= line_G05[32];	11'd426:G <= line_G05[22];	11'd436:G <= line_G05[12];	11'd446:G <= line_G05[2];
				11'd417:G <= line_G05[31];	11'd427:G <= line_G05[21];	11'd437:G <= line_G05[11];	11'd447:G <= line_G05[1];
				11'd418:G <= line_G05[30];	11'd428:G <= line_G05[20];	11'd438:G <= line_G05[10];	11'd448:G <= line_G05[0];
				default:G <= 0;
			endcase
		11'd328:
			case (pixel_col)
				11'd409:G <= line_G06[39];	11'd419:G <= line_G06[29];	11'd429:G <= line_G06[19];	11'd439:G <= line_G06[9];
				11'd410:G <= line_G06[38];	11'd420:G <= line_G06[28];	11'd430:G <= line_G06[18];	11'd440:G <= line_G06[8];
				11'd411:G <= line_G06[37];	11'd421:G <= line_G06[27];	11'd431:G <= line_G06[17];	11'd441:G <= line_G06[7];
				11'd412:G <= line_G06[36];	11'd422:G <= line_G06[26];	11'd432:G <= line_G06[16];	11'd442:G <= line_G06[6];
				11'd413:G <= line_G06[35];	11'd423:G <= line_G06[25];	11'd433:G <= line_G06[15];	11'd443:G <= line_G06[5];
				11'd414:G <= line_G06[34];	11'd424:G <= line_G06[24];	11'd434:G <= line_G06[14];	11'd444:G <= line_G06[4];
				11'd415:G <= line_G06[33];	11'd425:G <= line_G06[23];	11'd435:G <= line_G06[13];	11'd445:G <= line_G06[3];
				11'd416:G <= line_G06[32];	11'd426:G <= line_G06[22];	11'd436:G <= line_G06[12];	11'd446:G <= line_G06[2];
				11'd417:G <= line_G06[31];	11'd427:G <= line_G06[21];	11'd437:G <= line_G06[11];	11'd447:G <= line_G06[1];
				11'd418:G <= line_G06[30];	11'd428:G <= line_G06[20];	11'd438:G <= line_G06[10];	11'd448:G <= line_G06[0];
				default:G <= 0;
			endcase
		11'd329:
			case (pixel_col)
				11'd409:G <= line_G07[39];	11'd419:G <= line_G07[29];	11'd429:G <= line_G07[19];	11'd439:G <= line_G07[9];
				11'd410:G <= line_G07[38];	11'd420:G <= line_G07[28];	11'd430:G <= line_G07[18];	11'd440:G <= line_G07[8];
				11'd411:G <= line_G07[37];	11'd421:G <= line_G07[27];	11'd431:G <= line_G07[17];	11'd441:G <= line_G07[7];
				11'd412:G <= line_G07[36];	11'd422:G <= line_G07[26];	11'd432:G <= line_G07[16];	11'd442:G <= line_G07[6];
				11'd413:G <= line_G07[35];	11'd423:G <= line_G07[25];	11'd433:G <= line_G07[15];	11'd443:G <= line_G07[5];
				11'd414:G <= line_G07[34];	11'd424:G <= line_G07[24];	11'd434:G <= line_G07[14];	11'd444:G <= line_G07[4];
				11'd415:G <= line_G07[33];	11'd425:G <= line_G07[23];	11'd435:G <= line_G07[13];	11'd445:G <= line_G07[3];
				11'd416:G <= line_G07[32];	11'd426:G <= line_G07[22];	11'd436:G <= line_G07[12];	11'd446:G <= line_G07[2];
				11'd417:G <= line_G07[31];	11'd427:G <= line_G07[21];	11'd437:G <= line_G07[11];	11'd447:G <= line_G07[1];
				11'd418:G <= line_G07[30];	11'd428:G <= line_G07[20];	11'd438:G <= line_G07[10];	11'd448:G <= line_G07[0];
				default:G <= 0;
			endcase
		11'd330:
			case (pixel_col)
				11'd409:G <= line_G08[39];	11'd419:G <= line_G08[29];	11'd429:G <= line_G08[19];	11'd439:G <= line_G08[9];
				11'd410:G <= line_G08[38];	11'd420:G <= line_G08[28];	11'd430:G <= line_G08[18];	11'd440:G <= line_G08[8];
				11'd411:G <= line_G08[37];	11'd421:G <= line_G08[27];	11'd431:G <= line_G08[17];	11'd441:G <= line_G08[7];
				11'd412:G <= line_G08[36];	11'd422:G <= line_G08[26];	11'd432:G <= line_G08[16];	11'd442:G <= line_G08[6];
				11'd413:G <= line_G08[35];	11'd423:G <= line_G08[25];	11'd433:G <= line_G08[15];	11'd443:G <= line_G08[5];
				11'd414:G <= line_G08[34];	11'd424:G <= line_G08[24];	11'd434:G <= line_G08[14];	11'd444:G <= line_G08[4];
				11'd415:G <= line_G08[33];	11'd425:G <= line_G08[23];	11'd435:G <= line_G08[13];	11'd445:G <= line_G08[3];
				11'd416:G <= line_G08[32];	11'd426:G <= line_G08[22];	11'd436:G <= line_G08[12];	11'd446:G <= line_G08[2];
				11'd417:G <= line_G08[31];	11'd427:G <= line_G08[21];	11'd437:G <= line_G08[11];	11'd447:G <= line_G08[1];
				11'd418:G <= line_G08[30];	11'd428:G <= line_G08[20];	11'd438:G <= line_G08[10];	11'd448:G <= line_G08[0];
				default:G <= 0;
			endcase
		11'd331:
			case (pixel_col)
				11'd409:G <= line_G09[39];	11'd419:G <= line_G09[29];	11'd429:G <= line_G09[19];	11'd439:G <= line_G09[9];
				11'd410:G <= line_G09[38];	11'd420:G <= line_G09[28];	11'd430:G <= line_G09[18];	11'd440:G <= line_G09[8];
				11'd411:G <= line_G09[37];	11'd421:G <= line_G09[27];	11'd431:G <= line_G09[17];	11'd441:G <= line_G09[7];
				11'd412:G <= line_G09[36];	11'd422:G <= line_G09[26];	11'd432:G <= line_G09[16];	11'd442:G <= line_G09[6];
				11'd413:G <= line_G09[35];	11'd423:G <= line_G09[25];	11'd433:G <= line_G09[15];	11'd443:G <= line_G09[5];
				11'd414:G <= line_G09[34];	11'd424:G <= line_G09[24];	11'd434:G <= line_G09[14];	11'd444:G <= line_G09[4];
				11'd415:G <= line_G09[33];	11'd425:G <= line_G09[23];	11'd435:G <= line_G09[13];	11'd445:G <= line_G09[3];
				11'd416:G <= line_G09[32];	11'd426:G <= line_G09[22];	11'd436:G <= line_G09[12];	11'd446:G <= line_G09[2];
				11'd417:G <= line_G09[31];	11'd427:G <= line_G09[21];	11'd437:G <= line_G09[11];	11'd447:G <= line_G09[1];
				11'd418:G <= line_G09[30];	11'd428:G <= line_G09[20];	11'd438:G <= line_G09[10];	11'd448:G <= line_G09[0];
				default:G <= 0;
			endcase
		11'd332:
			case (pixel_col)
				11'd409:G <= line_G10[39];	11'd419:G <= line_G10[29];	11'd429:G <= line_G10[19];	11'd439:G <= line_G10[9];
				11'd410:G <= line_G10[38];	11'd420:G <= line_G10[28];	11'd430:G <= line_G10[18];	11'd440:G <= line_G10[8];
				11'd411:G <= line_G10[37];	11'd421:G <= line_G10[27];	11'd431:G <= line_G10[17];	11'd441:G <= line_G10[7];
				11'd412:G <= line_G10[36];	11'd422:G <= line_G10[26];	11'd432:G <= line_G10[16];	11'd442:G <= line_G10[6];
				11'd413:G <= line_G10[35];	11'd423:G <= line_G10[25];	11'd433:G <= line_G10[15];	11'd443:G <= line_G10[5];
				11'd414:G <= line_G10[34];	11'd424:G <= line_G10[24];	11'd434:G <= line_G10[14];	11'd444:G <= line_G10[4];
				11'd415:G <= line_G10[33];	11'd425:G <= line_G10[23];	11'd435:G <= line_G10[13];	11'd445:G <= line_G10[3];
				11'd416:G <= line_G10[32];	11'd426:G <= line_G10[22];	11'd436:G <= line_G10[12];	11'd446:G <= line_G10[2];
				11'd417:G <= line_G10[31];	11'd427:G <= line_G10[21];	11'd437:G <= line_G10[11];	11'd447:G <= line_G10[1];
				11'd418:G <= line_G10[30];	11'd428:G <= line_G10[20];	11'd438:G <= line_G10[10];	11'd448:G <= line_G10[0];
				default:G <= 0;
			endcase
		11'd333:
			case (pixel_col)
				11'd409:G <= line_G11[39];	11'd419:G <= line_G11[29];	11'd429:G <= line_G11[19];	11'd439:G <= line_G11[9];
				11'd410:G <= line_G11[38];	11'd420:G <= line_G11[28];	11'd430:G <= line_G11[18];	11'd440:G <= line_G11[8];
				11'd411:G <= line_G11[37];	11'd421:G <= line_G11[27];	11'd431:G <= line_G11[17];	11'd441:G <= line_G11[7];
				11'd412:G <= line_G11[36];	11'd422:G <= line_G11[26];	11'd432:G <= line_G11[16];	11'd442:G <= line_G11[6];
				11'd413:G <= line_G11[35];	11'd423:G <= line_G11[25];	11'd433:G <= line_G11[15];	11'd443:G <= line_G11[5];
				11'd414:G <= line_G11[34];	11'd424:G <= line_G11[24];	11'd434:G <= line_G11[14];	11'd444:G <= line_G11[4];
				11'd415:G <= line_G11[33];	11'd425:G <= line_G11[23];	11'd435:G <= line_G11[13];	11'd445:G <= line_G11[3];
				11'd416:G <= line_G11[32];	11'd426:G <= line_G11[22];	11'd436:G <= line_G11[12];	11'd446:G <= line_G11[2];
				11'd417:G <= line_G11[31];	11'd427:G <= line_G11[21];	11'd437:G <= line_G11[11];	11'd447:G <= line_G11[1];
				11'd418:G <= line_G11[30];	11'd428:G <= line_G11[20];	11'd438:G <= line_G11[10];	11'd448:G <= line_G11[0];
				default:G <= 0;
			endcase
		11'd334:
			case (pixel_col)
				11'd409:G <= line_G12[39];	11'd419:G <= line_G12[29];	11'd429:G <= line_G12[19];	11'd439:G <= line_G12[9];
				11'd410:G <= line_G12[38];	11'd420:G <= line_G12[28];	11'd430:G <= line_G12[18];	11'd440:G <= line_G12[8];
				11'd411:G <= line_G12[37];	11'd421:G <= line_G12[27];	11'd431:G <= line_G12[17];	11'd441:G <= line_G12[7];
				11'd412:G <= line_G12[36];	11'd422:G <= line_G12[26];	11'd432:G <= line_G12[16];	11'd442:G <= line_G12[6];
				11'd413:G <= line_G12[35];	11'd423:G <= line_G12[25];	11'd433:G <= line_G12[15];	11'd443:G <= line_G12[5];
				11'd414:G <= line_G12[34];	11'd424:G <= line_G12[24];	11'd434:G <= line_G12[14];	11'd444:G <= line_G12[4];
				11'd415:G <= line_G12[33];	11'd425:G <= line_G12[23];	11'd435:G <= line_G12[13];	11'd445:G <= line_G12[3];
				11'd416:G <= line_G12[32];	11'd426:G <= line_G12[22];	11'd436:G <= line_G12[12];	11'd446:G <= line_G12[2];
				11'd417:G <= line_G12[31];	11'd427:G <= line_G12[21];	11'd437:G <= line_G12[11];	11'd447:G <= line_G12[1];
				11'd418:G <= line_G12[30];	11'd428:G <= line_G12[20];	11'd438:G <= line_G12[10];	11'd448:G <= line_G12[0];
				default:G <= 0;
			endcase
		11'd335:
			case (pixel_col)
				11'd409:G <= line_G13[39];	11'd419:G <= line_G13[29];	11'd429:G <= line_G13[19];	11'd439:G <= line_G13[9];
				11'd410:G <= line_G13[38];	11'd420:G <= line_G13[28];	11'd430:G <= line_G13[18];	11'd440:G <= line_G13[8];
				11'd411:G <= line_G13[37];	11'd421:G <= line_G13[27];	11'd431:G <= line_G13[17];	11'd441:G <= line_G13[7];
				11'd412:G <= line_G13[36];	11'd422:G <= line_G13[26];	11'd432:G <= line_G13[16];	11'd442:G <= line_G13[6];
				11'd413:G <= line_G13[35];	11'd423:G <= line_G13[25];	11'd433:G <= line_G13[15];	11'd443:G <= line_G13[5];
				11'd414:G <= line_G13[34];	11'd424:G <= line_G13[24];	11'd434:G <= line_G13[14];	11'd444:G <= line_G13[4];
				11'd415:G <= line_G13[33];	11'd425:G <= line_G13[23];	11'd435:G <= line_G13[13];	11'd445:G <= line_G13[3];
				11'd416:G <= line_G13[32];	11'd426:G <= line_G13[22];	11'd436:G <= line_G13[12];	11'd446:G <= line_G13[2];
				11'd417:G <= line_G13[31];	11'd427:G <= line_G13[21];	11'd437:G <= line_G13[11];	11'd447:G <= line_G13[1];
				11'd418:G <= line_G13[30];	11'd428:G <= line_G13[20];	11'd438:G <= line_G13[10];	11'd448:G <= line_G13[0];
				default:G <= 0;
			endcase
		11'd336:
			case (pixel_col)
				11'd409:G <= line_G14[39];	11'd419:G <= line_G14[29];	11'd429:G <= line_G14[19];	11'd439:G <= line_G14[9];
				11'd410:G <= line_G14[38];	11'd420:G <= line_G14[28];	11'd430:G <= line_G14[18];	11'd440:G <= line_G14[8];
				11'd411:G <= line_G14[37];	11'd421:G <= line_G14[27];	11'd431:G <= line_G14[17];	11'd441:G <= line_G14[7];
				11'd412:G <= line_G14[36];	11'd422:G <= line_G14[26];	11'd432:G <= line_G14[16];	11'd442:G <= line_G14[6];
				11'd413:G <= line_G14[35];	11'd423:G <= line_G14[25];	11'd433:G <= line_G14[15];	11'd443:G <= line_G14[5];
				11'd414:G <= line_G14[34];	11'd424:G <= line_G14[24];	11'd434:G <= line_G14[14];	11'd444:G <= line_G14[4];
				11'd415:G <= line_G14[33];	11'd425:G <= line_G14[23];	11'd435:G <= line_G14[13];	11'd445:G <= line_G14[3];
				11'd416:G <= line_G14[32];	11'd426:G <= line_G14[22];	11'd436:G <= line_G14[12];	11'd446:G <= line_G14[2];
				11'd417:G <= line_G14[31];	11'd427:G <= line_G14[21];	11'd437:G <= line_G14[11];	11'd447:G <= line_G14[1];
				11'd418:G <= line_G14[30];	11'd428:G <= line_G14[20];	11'd438:G <= line_G14[10];	11'd448:G <= line_G14[0];
				default:G <= 0;
			endcase
		11'd337:
			case (pixel_col)
				11'd409:G <= line_G15[39];	11'd419:G <= line_G15[29];	11'd429:G <= line_G15[19];	11'd439:G <= line_G15[9];
				11'd410:G <= line_G15[38];	11'd420:G <= line_G15[28];	11'd430:G <= line_G15[18];	11'd440:G <= line_G15[8];
				11'd411:G <= line_G15[37];	11'd421:G <= line_G15[27];	11'd431:G <= line_G15[17];	11'd441:G <= line_G15[7];
				11'd412:G <= line_G15[36];	11'd422:G <= line_G15[26];	11'd432:G <= line_G15[16];	11'd442:G <= line_G15[6];
				11'd413:G <= line_G15[35];	11'd423:G <= line_G15[25];	11'd433:G <= line_G15[15];	11'd443:G <= line_G15[5];
				11'd414:G <= line_G15[34];	11'd424:G <= line_G15[24];	11'd434:G <= line_G15[14];	11'd444:G <= line_G15[4];
				11'd415:G <= line_G15[33];	11'd425:G <= line_G15[23];	11'd435:G <= line_G15[13];	11'd445:G <= line_G15[3];
				11'd416:G <= line_G15[32];	11'd426:G <= line_G15[22];	11'd436:G <= line_G15[12];	11'd446:G <= line_G15[2];
				11'd417:G <= line_G15[31];	11'd427:G <= line_G15[21];	11'd437:G <= line_G15[11];	11'd447:G <= line_G15[1];
				11'd418:G <= line_G15[30];	11'd428:G <= line_G15[20];	11'd438:G <= line_G15[10];	11'd448:G <= line_G15[0];
				default:G <= 0;
			endcase
		default:G <= 0;
	endcase
end


always @(posedge clk) begin
	case (pixel_row)
		11'd323:
			case (pixel_col)
				11'd459:A <= line_A01[39];	11'd469:A <= line_A01[29];	11'd479:A <= line_A01[19];	11'd489:A <= line_A01[9];
				11'd460:A <= line_A01[38];	11'd470:A <= line_A01[28];	11'd480:A <= line_A01[18];	11'd490:A <= line_A01[8];
				11'd461:A <= line_A01[37];	11'd471:A <= line_A01[27];	11'd481:A <= line_A01[17];	11'd491:A <= line_A01[7];
				11'd462:A <= line_A01[36];	11'd472:A <= line_A01[26];	11'd482:A <= line_A01[16];	11'd492:A <= line_A01[6];
				11'd463:A <= line_A01[35];	11'd473:A <= line_A01[25];	11'd483:A <= line_A01[15];	11'd493:A <= line_A01[5];
				11'd464:A <= line_A01[34];	11'd474:A <= line_A01[24];	11'd484:A <= line_A01[14];	11'd494:A <= line_A01[4];
				11'd465:A <= line_A01[33];	11'd475:A <= line_A01[23];	11'd485:A <= line_A01[13];	11'd495:A <= line_A01[3];
				11'd466:A <= line_A01[32];	11'd476:A <= line_A01[22];	11'd486:A <= line_A01[12];	11'd496:A <= line_A01[2];
				11'd467:A <= line_A01[31];	11'd477:A <= line_A01[21];	11'd487:A <= line_A01[11];	11'd497:A <= line_A01[1];
				11'd468:A <= line_A01[30];	11'd478:A <= line_A01[20];	11'd488:A <= line_A01[10];	11'd498:A <= line_A01[0];
				default:A <= 0;
			endcase
		11'd324:
			case (pixel_col)
				11'd459:A <= line_A02[39];	11'd469:A <= line_A02[29];	11'd479:A <= line_A02[19];	11'd489:A <= line_A02[9];
				11'd460:A <= line_A02[38];	11'd470:A <= line_A02[28];	11'd480:A <= line_A02[18];	11'd490:A <= line_A02[8];
				11'd461:A <= line_A02[37];	11'd471:A <= line_A02[27];	11'd481:A <= line_A02[17];	11'd491:A <= line_A02[7];
				11'd462:A <= line_A02[36];	11'd472:A <= line_A02[26];	11'd482:A <= line_A02[16];	11'd492:A <= line_A02[6];
				11'd463:A <= line_A02[35];	11'd473:A <= line_A02[25];	11'd483:A <= line_A02[15];	11'd493:A <= line_A02[5];
				11'd464:A <= line_A02[34];	11'd474:A <= line_A02[24];	11'd484:A <= line_A02[14];	11'd494:A <= line_A02[4];
				11'd465:A <= line_A02[33];	11'd475:A <= line_A02[23];	11'd485:A <= line_A02[13];	11'd495:A <= line_A02[3];
				11'd466:A <= line_A02[32];	11'd476:A <= line_A02[22];	11'd486:A <= line_A02[12];	11'd496:A <= line_A02[2];
				11'd467:A <= line_A02[31];	11'd477:A <= line_A02[21];	11'd487:A <= line_A02[11];	11'd497:A <= line_A02[1];
				11'd468:A <= line_A02[30];	11'd478:A <= line_A02[20];	11'd488:A <= line_A02[10];	11'd498:A <= line_A02[0];
				default:A <= 0;
			endcase
		11'd325:
			case (pixel_col)
				11'd459:A <= line_A03[39];	11'd469:A <= line_A03[29];	11'd479:A <= line_A03[19];	11'd489:A <= line_A03[9];
				11'd460:A <= line_A03[38];	11'd470:A <= line_A03[28];	11'd480:A <= line_A03[18];	11'd490:A <= line_A03[8];
				11'd461:A <= line_A03[37];	11'd471:A <= line_A03[27];	11'd481:A <= line_A03[17];	11'd491:A <= line_A03[7];
				11'd462:A <= line_A03[36];	11'd472:A <= line_A03[26];	11'd482:A <= line_A03[16];	11'd492:A <= line_A03[6];
				11'd463:A <= line_A03[35];	11'd473:A <= line_A03[25];	11'd483:A <= line_A03[15];	11'd493:A <= line_A03[5];
				11'd464:A <= line_A03[34];	11'd474:A <= line_A03[24];	11'd484:A <= line_A03[14];	11'd494:A <= line_A03[4];
				11'd465:A <= line_A03[33];	11'd475:A <= line_A03[23];	11'd485:A <= line_A03[13];	11'd495:A <= line_A03[3];
				11'd466:A <= line_A03[32];	11'd476:A <= line_A03[22];	11'd486:A <= line_A03[12];	11'd496:A <= line_A03[2];
				11'd467:A <= line_A03[31];	11'd477:A <= line_A03[21];	11'd487:A <= line_A03[11];	11'd497:A <= line_A03[1];
				11'd468:A <= line_A03[30];	11'd478:A <= line_A03[20];	11'd488:A <= line_A03[10];	11'd498:A <= line_A03[0];
				default:A <= 0;
			endcase
		11'd326:
			case (pixel_col)
				11'd459:A <= line_A04[39];	11'd469:A <= line_A04[29];	11'd479:A <= line_A04[19];	11'd489:A <= line_A04[9];
				11'd460:A <= line_A04[38];	11'd470:A <= line_A04[28];	11'd480:A <= line_A04[18];	11'd490:A <= line_A04[8];
				11'd461:A <= line_A04[37];	11'd471:A <= line_A04[27];	11'd481:A <= line_A04[17];	11'd491:A <= line_A04[7];
				11'd462:A <= line_A04[36];	11'd472:A <= line_A04[26];	11'd482:A <= line_A04[16];	11'd492:A <= line_A04[6];
				11'd463:A <= line_A04[35];	11'd473:A <= line_A04[25];	11'd483:A <= line_A04[15];	11'd493:A <= line_A04[5];
				11'd464:A <= line_A04[34];	11'd474:A <= line_A04[24];	11'd484:A <= line_A04[14];	11'd494:A <= line_A04[4];
				11'd465:A <= line_A04[33];	11'd475:A <= line_A04[23];	11'd485:A <= line_A04[13];	11'd495:A <= line_A04[3];
				11'd466:A <= line_A04[32];	11'd476:A <= line_A04[22];	11'd486:A <= line_A04[12];	11'd496:A <= line_A04[2];
				11'd467:A <= line_A04[31];	11'd477:A <= line_A04[21];	11'd487:A <= line_A04[11];	11'd497:A <= line_A04[1];
				11'd468:A <= line_A04[30];	11'd478:A <= line_A04[20];	11'd488:A <= line_A04[10];	11'd498:A <= line_A04[0];
				default:A <= 0;
			endcase
		11'd327:
			case (pixel_col)
				11'd459:A <= line_A05[39];	11'd469:A <= line_A05[29];	11'd479:A <= line_A05[19];	11'd489:A <= line_A05[9];
				11'd460:A <= line_A05[38];	11'd470:A <= line_A05[28];	11'd480:A <= line_A05[18];	11'd490:A <= line_A05[8];
				11'd461:A <= line_A05[37];	11'd471:A <= line_A05[27];	11'd481:A <= line_A05[17];	11'd491:A <= line_A05[7];
				11'd462:A <= line_A05[36];	11'd472:A <= line_A05[26];	11'd482:A <= line_A05[16];	11'd492:A <= line_A05[6];
				11'd463:A <= line_A05[35];	11'd473:A <= line_A05[25];	11'd483:A <= line_A05[15];	11'd493:A <= line_A05[5];
				11'd464:A <= line_A05[34];	11'd474:A <= line_A05[24];	11'd484:A <= line_A05[14];	11'd494:A <= line_A05[4];
				11'd465:A <= line_A05[33];	11'd475:A <= line_A05[23];	11'd485:A <= line_A05[13];	11'd495:A <= line_A05[3];
				11'd466:A <= line_A05[32];	11'd476:A <= line_A05[22];	11'd486:A <= line_A05[12];	11'd496:A <= line_A05[2];
				11'd467:A <= line_A05[31];	11'd477:A <= line_A05[21];	11'd487:A <= line_A05[11];	11'd497:A <= line_A05[1];
				11'd468:A <= line_A05[30];	11'd478:A <= line_A05[20];	11'd488:A <= line_A05[10];	11'd498:A <= line_A05[0];
				default:A <= 0;
			endcase
		11'd328:
			case (pixel_col)
				11'd459:A <= line_A06[39];	11'd469:A <= line_A06[29];	11'd479:A <= line_A06[19];	11'd489:A <= line_A06[9];
				11'd460:A <= line_A06[38];	11'd470:A <= line_A06[28];	11'd480:A <= line_A06[18];	11'd490:A <= line_A06[8];
				11'd461:A <= line_A06[37];	11'd471:A <= line_A06[27];	11'd481:A <= line_A06[17];	11'd491:A <= line_A06[7];
				11'd462:A <= line_A06[36];	11'd472:A <= line_A06[26];	11'd482:A <= line_A06[16];	11'd492:A <= line_A06[6];
				11'd463:A <= line_A06[35];	11'd473:A <= line_A06[25];	11'd483:A <= line_A06[15];	11'd493:A <= line_A06[5];
				11'd464:A <= line_A06[34];	11'd474:A <= line_A06[24];	11'd484:A <= line_A06[14];	11'd494:A <= line_A06[4];
				11'd465:A <= line_A06[33];	11'd475:A <= line_A06[23];	11'd485:A <= line_A06[13];	11'd495:A <= line_A06[3];
				11'd466:A <= line_A06[32];	11'd476:A <= line_A06[22];	11'd486:A <= line_A06[12];	11'd496:A <= line_A06[2];
				11'd467:A <= line_A06[31];	11'd477:A <= line_A06[21];	11'd487:A <= line_A06[11];	11'd497:A <= line_A06[1];
				11'd468:A <= line_A06[30];	11'd478:A <= line_A06[20];	11'd488:A <= line_A06[10];	11'd498:A <= line_A06[0];
				default:A <= 0;
			endcase
		11'd329:
			case (pixel_col)
				11'd459:A <= line_A07[39];	11'd469:A <= line_A07[29];	11'd479:A <= line_A07[19];	11'd489:A <= line_A07[9];
				11'd460:A <= line_A07[38];	11'd470:A <= line_A07[28];	11'd480:A <= line_A07[18];	11'd490:A <= line_A07[8];
				11'd461:A <= line_A07[37];	11'd471:A <= line_A07[27];	11'd481:A <= line_A07[17];	11'd491:A <= line_A07[7];
				11'd462:A <= line_A07[36];	11'd472:A <= line_A07[26];	11'd482:A <= line_A07[16];	11'd492:A <= line_A07[6];
				11'd463:A <= line_A07[35];	11'd473:A <= line_A07[25];	11'd483:A <= line_A07[15];	11'd493:A <= line_A07[5];
				11'd464:A <= line_A07[34];	11'd474:A <= line_A07[24];	11'd484:A <= line_A07[14];	11'd494:A <= line_A07[4];
				11'd465:A <= line_A07[33];	11'd475:A <= line_A07[23];	11'd485:A <= line_A07[13];	11'd495:A <= line_A07[3];
				11'd466:A <= line_A07[32];	11'd476:A <= line_A07[22];	11'd486:A <= line_A07[12];	11'd496:A <= line_A07[2];
				11'd467:A <= line_A07[31];	11'd477:A <= line_A07[21];	11'd487:A <= line_A07[11];	11'd497:A <= line_A07[1];
				11'd468:A <= line_A07[30];	11'd478:A <= line_A07[20];	11'd488:A <= line_A07[10];	11'd498:A <= line_A07[0];
				default:A <= 0;
			endcase
		11'd330:
			case (pixel_col)
				11'd459:A <= line_A08[39];	11'd469:A <= line_A08[29];	11'd479:A <= line_A08[19];	11'd489:A <= line_A08[9];
				11'd460:A <= line_A08[38];	11'd470:A <= line_A08[28];	11'd480:A <= line_A08[18];	11'd490:A <= line_A08[8];
				11'd461:A <= line_A08[37];	11'd471:A <= line_A08[27];	11'd481:A <= line_A08[17];	11'd491:A <= line_A08[7];
				11'd462:A <= line_A08[36];	11'd472:A <= line_A08[26];	11'd482:A <= line_A08[16];	11'd492:A <= line_A08[6];
				11'd463:A <= line_A08[35];	11'd473:A <= line_A08[25];	11'd483:A <= line_A08[15];	11'd493:A <= line_A08[5];
				11'd464:A <= line_A08[34];	11'd474:A <= line_A08[24];	11'd484:A <= line_A08[14];	11'd494:A <= line_A08[4];
				11'd465:A <= line_A08[33];	11'd475:A <= line_A08[23];	11'd485:A <= line_A08[13];	11'd495:A <= line_A08[3];
				11'd466:A <= line_A08[32];	11'd476:A <= line_A08[22];	11'd486:A <= line_A08[12];	11'd496:A <= line_A08[2];
				11'd467:A <= line_A08[31];	11'd477:A <= line_A08[21];	11'd487:A <= line_A08[11];	11'd497:A <= line_A08[1];
				11'd468:A <= line_A08[30];	11'd478:A <= line_A08[20];	11'd488:A <= line_A08[10];	11'd498:A <= line_A08[0];
				default:A <= 0;
			endcase
		11'd331:
			case (pixel_col)
				11'd459:A <= line_A09[39];	11'd469:A <= line_A09[29];	11'd479:A <= line_A09[19];	11'd489:A <= line_A09[9];
				11'd460:A <= line_A09[38];	11'd470:A <= line_A09[28];	11'd480:A <= line_A09[18];	11'd490:A <= line_A09[8];
				11'd461:A <= line_A09[37];	11'd471:A <= line_A09[27];	11'd481:A <= line_A09[17];	11'd491:A <= line_A09[7];
				11'd462:A <= line_A09[36];	11'd472:A <= line_A09[26];	11'd482:A <= line_A09[16];	11'd492:A <= line_A09[6];
				11'd463:A <= line_A09[35];	11'd473:A <= line_A09[25];	11'd483:A <= line_A09[15];	11'd493:A <= line_A09[5];
				11'd464:A <= line_A09[34];	11'd474:A <= line_A09[24];	11'd484:A <= line_A09[14];	11'd494:A <= line_A09[4];
				11'd465:A <= line_A09[33];	11'd475:A <= line_A09[23];	11'd485:A <= line_A09[13];	11'd495:A <= line_A09[3];
				11'd466:A <= line_A09[32];	11'd476:A <= line_A09[22];	11'd486:A <= line_A09[12];	11'd496:A <= line_A09[2];
				11'd467:A <= line_A09[31];	11'd477:A <= line_A09[21];	11'd487:A <= line_A09[11];	11'd497:A <= line_A09[1];
				11'd468:A <= line_A09[30];	11'd478:A <= line_A09[20];	11'd488:A <= line_A09[10];	11'd498:A <= line_A09[0];
				default:A <= 0;
			endcase
		11'd332:
			case (pixel_col)
				11'd459:A <= line_A10[39];	11'd469:A <= line_A10[29];	11'd479:A <= line_A10[19];	11'd489:A <= line_A10[9];
				11'd460:A <= line_A10[38];	11'd470:A <= line_A10[28];	11'd480:A <= line_A10[18];	11'd490:A <= line_A10[8];
				11'd461:A <= line_A10[37];	11'd471:A <= line_A10[27];	11'd481:A <= line_A10[17];	11'd491:A <= line_A10[7];
				11'd462:A <= line_A10[36];	11'd472:A <= line_A10[26];	11'd482:A <= line_A10[16];	11'd492:A <= line_A10[6];
				11'd463:A <= line_A10[35];	11'd473:A <= line_A10[25];	11'd483:A <= line_A10[15];	11'd493:A <= line_A10[5];
				11'd464:A <= line_A10[34];	11'd474:A <= line_A10[24];	11'd484:A <= line_A10[14];	11'd494:A <= line_A10[4];
				11'd465:A <= line_A10[33];	11'd475:A <= line_A10[23];	11'd485:A <= line_A10[13];	11'd495:A <= line_A10[3];
				11'd466:A <= line_A10[32];	11'd476:A <= line_A10[22];	11'd486:A <= line_A10[12];	11'd496:A <= line_A10[2];
				11'd467:A <= line_A10[31];	11'd477:A <= line_A10[21];	11'd487:A <= line_A10[11];	11'd497:A <= line_A10[1];
				11'd468:A <= line_A10[30];	11'd478:A <= line_A10[20];	11'd488:A <= line_A10[10];	11'd498:A <= line_A10[0];
				default:A <= 0;
			endcase
		11'd333:
			case (pixel_col)
				11'd459:A <= line_A11[39];	11'd469:A <= line_A11[29];	11'd479:A <= line_A11[19];	11'd489:A <= line_A11[9];
				11'd460:A <= line_A11[38];	11'd470:A <= line_A11[28];	11'd480:A <= line_A11[18];	11'd490:A <= line_A11[8];
				11'd461:A <= line_A11[37];	11'd471:A <= line_A11[27];	11'd481:A <= line_A11[17];	11'd491:A <= line_A11[7];
				11'd462:A <= line_A11[36];	11'd472:A <= line_A11[26];	11'd482:A <= line_A11[16];	11'd492:A <= line_A11[6];
				11'd463:A <= line_A11[35];	11'd473:A <= line_A11[25];	11'd483:A <= line_A11[15];	11'd493:A <= line_A11[5];
				11'd464:A <= line_A11[34];	11'd474:A <= line_A11[24];	11'd484:A <= line_A11[14];	11'd494:A <= line_A11[4];
				11'd465:A <= line_A11[33];	11'd475:A <= line_A11[23];	11'd485:A <= line_A11[13];	11'd495:A <= line_A11[3];
				11'd466:A <= line_A11[32];	11'd476:A <= line_A11[22];	11'd486:A <= line_A11[12];	11'd496:A <= line_A11[2];
				11'd467:A <= line_A11[31];	11'd477:A <= line_A11[21];	11'd487:A <= line_A11[11];	11'd497:A <= line_A11[1];
				11'd468:A <= line_A11[30];	11'd478:A <= line_A11[20];	11'd488:A <= line_A11[10];	11'd498:A <= line_A11[0];
				default:A <= 0;
			endcase
		11'd334:
			case (pixel_col)
				11'd459:A <= line_A12[39];	11'd469:A <= line_A12[29];	11'd479:A <= line_A12[19];	11'd489:A <= line_A12[9];
				11'd460:A <= line_A12[38];	11'd470:A <= line_A12[28];	11'd480:A <= line_A12[18];	11'd490:A <= line_A12[8];
				11'd461:A <= line_A12[37];	11'd471:A <= line_A12[27];	11'd481:A <= line_A12[17];	11'd491:A <= line_A12[7];
				11'd462:A <= line_A12[36];	11'd472:A <= line_A12[26];	11'd482:A <= line_A12[16];	11'd492:A <= line_A12[6];
				11'd463:A <= line_A12[35];	11'd473:A <= line_A12[25];	11'd483:A <= line_A12[15];	11'd493:A <= line_A12[5];
				11'd464:A <= line_A12[34];	11'd474:A <= line_A12[24];	11'd484:A <= line_A12[14];	11'd494:A <= line_A12[4];
				11'd465:A <= line_A12[33];	11'd475:A <= line_A12[23];	11'd485:A <= line_A12[13];	11'd495:A <= line_A12[3];
				11'd466:A <= line_A12[32];	11'd476:A <= line_A12[22];	11'd486:A <= line_A12[12];	11'd496:A <= line_A12[2];
				11'd467:A <= line_A12[31];	11'd477:A <= line_A12[21];	11'd487:A <= line_A12[11];	11'd497:A <= line_A12[1];
				11'd468:A <= line_A12[30];	11'd478:A <= line_A12[20];	11'd488:A <= line_A12[10];	11'd498:A <= line_A12[0];
				default:A <= 0;
			endcase
		11'd335:
			case (pixel_col)
				11'd459:A <= line_A13[39];	11'd469:A <= line_A13[29];	11'd479:A <= line_A13[19];	11'd489:A <= line_A13[9];
				11'd460:A <= line_A13[38];	11'd470:A <= line_A13[28];	11'd480:A <= line_A13[18];	11'd490:A <= line_A13[8];
				11'd461:A <= line_A13[37];	11'd471:A <= line_A13[27];	11'd481:A <= line_A13[17];	11'd491:A <= line_A13[7];
				11'd462:A <= line_A13[36];	11'd472:A <= line_A13[26];	11'd482:A <= line_A13[16];	11'd492:A <= line_A13[6];
				11'd463:A <= line_A13[35];	11'd473:A <= line_A13[25];	11'd483:A <= line_A13[15];	11'd493:A <= line_A13[5];
				11'd464:A <= line_A13[34];	11'd474:A <= line_A13[24];	11'd484:A <= line_A13[14];	11'd494:A <= line_A13[4];
				11'd465:A <= line_A13[33];	11'd475:A <= line_A13[23];	11'd485:A <= line_A13[13];	11'd495:A <= line_A13[3];
				11'd466:A <= line_A13[32];	11'd476:A <= line_A13[22];	11'd486:A <= line_A13[12];	11'd496:A <= line_A13[2];
				11'd467:A <= line_A13[31];	11'd477:A <= line_A13[21];	11'd487:A <= line_A13[11];	11'd497:A <= line_A13[1];
				11'd468:A <= line_A13[30];	11'd478:A <= line_A13[20];	11'd488:A <= line_A13[10];	11'd498:A <= line_A13[0];
				default:A <= 0;
			endcase
		11'd336:
			case (pixel_col)
				11'd459:A <= line_A14[39];	11'd469:A <= line_A14[29];	11'd479:A <= line_A14[19];	11'd489:A <= line_A14[9];
				11'd460:A <= line_A14[38];	11'd470:A <= line_A14[28];	11'd480:A <= line_A14[18];	11'd490:A <= line_A14[8];
				11'd461:A <= line_A14[37];	11'd471:A <= line_A14[27];	11'd481:A <= line_A14[17];	11'd491:A <= line_A14[7];
				11'd462:A <= line_A14[36];	11'd472:A <= line_A14[26];	11'd482:A <= line_A14[16];	11'd492:A <= line_A14[6];
				11'd463:A <= line_A14[35];	11'd473:A <= line_A14[25];	11'd483:A <= line_A14[15];	11'd493:A <= line_A14[5];
				11'd464:A <= line_A14[34];	11'd474:A <= line_A14[24];	11'd484:A <= line_A14[14];	11'd494:A <= line_A14[4];
				11'd465:A <= line_A14[33];	11'd475:A <= line_A14[23];	11'd485:A <= line_A14[13];	11'd495:A <= line_A14[3];
				11'd466:A <= line_A14[32];	11'd476:A <= line_A14[22];	11'd486:A <= line_A14[12];	11'd496:A <= line_A14[2];
				11'd467:A <= line_A14[31];	11'd477:A <= line_A14[21];	11'd487:A <= line_A14[11];	11'd497:A <= line_A14[1];
				11'd468:A <= line_A14[30];	11'd478:A <= line_A14[20];	11'd488:A <= line_A14[10];	11'd498:A <= line_A14[0];
				default:A <= 0;
			endcase
		11'd337:
			case (pixel_col)
				11'd459:A <= line_A15[39];	11'd469:A <= line_A15[29];	11'd479:A <= line_A15[19];	11'd489:A <= line_A15[9];
				11'd460:A <= line_A15[38];	11'd470:A <= line_A15[28];	11'd480:A <= line_A15[18];	11'd490:A <= line_A15[8];
				11'd461:A <= line_A15[37];	11'd471:A <= line_A15[27];	11'd481:A <= line_A15[17];	11'd491:A <= line_A15[7];
				11'd462:A <= line_A15[36];	11'd472:A <= line_A15[26];	11'd482:A <= line_A15[16];	11'd492:A <= line_A15[6];
				11'd463:A <= line_A15[35];	11'd473:A <= line_A15[25];	11'd483:A <= line_A15[15];	11'd493:A <= line_A15[5];
				11'd464:A <= line_A15[34];	11'd474:A <= line_A15[24];	11'd484:A <= line_A15[14];	11'd494:A <= line_A15[4];
				11'd465:A <= line_A15[33];	11'd475:A <= line_A15[23];	11'd485:A <= line_A15[13];	11'd495:A <= line_A15[3];
				11'd466:A <= line_A15[32];	11'd476:A <= line_A15[22];	11'd486:A <= line_A15[12];	11'd496:A <= line_A15[2];
				11'd467:A <= line_A15[31];	11'd477:A <= line_A15[21];	11'd487:A <= line_A15[11];	11'd497:A <= line_A15[1];
				11'd468:A <= line_A15[30];	11'd478:A <= line_A15[20];	11'd488:A <= line_A15[10];	11'd498:A <= line_A15[0];
				default:A <= 0;
			endcase
		default:A <= 0;
	endcase
end


always @(posedge clk) begin

		case (pixel_row)
		11'd323:
			case (pixel_col)
				11'd509:M <= line_M01[39];	11'd519:M <= line_M01[29];	11'd529:M <= line_M01[19];	11'd539:M <= line_M01[9];
				11'd510:M <= line_M01[38];	11'd520:M <= line_M01[28];	11'd530:M <= line_M01[18];	11'd540:M <= line_M01[8];
				11'd511:M <= line_M01[37];	11'd521:M <= line_M01[27];	11'd531:M <= line_M01[17];	11'd541:M <= line_M01[7];
				11'd512:M <= line_M01[36];	11'd522:M <= line_M01[26];	11'd532:M <= line_M01[16];	11'd542:M <= line_M01[6];
				11'd513:M <= line_M01[35];	11'd523:M <= line_M01[25];	11'd533:M <= line_M01[15];	11'd543:M <= line_M01[5];
				11'd514:M <= line_M01[34];	11'd524:M <= line_M01[24];	11'd534:M <= line_M01[14];	11'd544:M <= line_M01[4];
				11'd515:M <= line_M01[33];	11'd525:M <= line_M01[23];	11'd535:M <= line_M01[13];	11'd545:M <= line_M01[3];
				11'd516:M <= line_M01[32];	11'd526:M <= line_M01[22];	11'd536:M <= line_M01[12];	11'd546:M <= line_M01[2];
				11'd517:M <= line_M01[31];	11'd527:M <= line_M01[21];	11'd537:M <= line_M01[11];	11'd547:M <= line_M01[1];
				11'd518:M <= line_M01[30];	11'd528:M <= line_M01[20];	11'd538:M <= line_M01[10];	11'd548:M <= line_M01[0];
				default:M <= 0;
			endcase
		11'd324:
			case (pixel_col)
				11'd509:M <= line_M02[39];	11'd519:M <= line_M02[29];	11'd529:M <= line_M02[19];	11'd539:M <= line_M02[9];
				11'd510:M <= line_M02[38];	11'd520:M <= line_M02[28];	11'd530:M <= line_M02[18];	11'd540:M <= line_M02[8];
				11'd511:M <= line_M02[37];	11'd521:M <= line_M02[27];	11'd531:M <= line_M02[17];	11'd541:M <= line_M02[7];
				11'd512:M <= line_M02[36];	11'd522:M <= line_M02[26];	11'd532:M <= line_M02[16];	11'd542:M <= line_M02[6];
				11'd513:M <= line_M02[35];	11'd523:M <= line_M02[25];	11'd533:M <= line_M02[15];	11'd543:M <= line_M02[5];
				11'd514:M <= line_M02[34];	11'd524:M <= line_M02[24];	11'd534:M <= line_M02[14];	11'd544:M <= line_M02[4];
				11'd515:M <= line_M02[33];	11'd525:M <= line_M02[23];	11'd535:M <= line_M02[13];	11'd545:M <= line_M02[3];
				11'd516:M <= line_M02[32];	11'd526:M <= line_M02[22];	11'd536:M <= line_M02[12];	11'd546:M <= line_M02[2];
				11'd517:M <= line_M02[31];	11'd527:M <= line_M02[21];	11'd537:M <= line_M02[11];	11'd547:M <= line_M02[1];
				11'd518:M <= line_M02[30];	11'd528:M <= line_M02[20];	11'd538:M <= line_M02[10];	11'd548:M <= line_M02[0];
				default:M <= 0;
			endcase
		11'd325:
			case (pixel_col)
				11'd509:M <= line_M03[39];	11'd519:M <= line_M03[29];	11'd529:M <= line_M03[19];	11'd539:M <= line_M03[9];
				11'd510:M <= line_M03[38];	11'd520:M <= line_M03[28];	11'd530:M <= line_M03[18];	11'd540:M <= line_M03[8];
				11'd511:M <= line_M03[37];	11'd521:M <= line_M03[27];	11'd531:M <= line_M03[17];	11'd541:M <= line_M03[7];
				11'd512:M <= line_M03[36];	11'd522:M <= line_M03[26];	11'd532:M <= line_M03[16];	11'd542:M <= line_M03[6];
				11'd513:M <= line_M03[35];	11'd523:M <= line_M03[25];	11'd533:M <= line_M03[15];	11'd543:M <= line_M03[5];
				11'd514:M <= line_M03[34];	11'd524:M <= line_M03[24];	11'd534:M <= line_M03[14];	11'd544:M <= line_M03[4];
				11'd515:M <= line_M03[33];	11'd525:M <= line_M03[23];	11'd535:M <= line_M03[13];	11'd545:M <= line_M03[3];
				11'd516:M <= line_M03[32];	11'd526:M <= line_M03[22];	11'd536:M <= line_M03[12];	11'd546:M <= line_M03[2];
				11'd517:M <= line_M03[31];	11'd527:M <= line_M03[21];	11'd537:M <= line_M03[11];	11'd547:M <= line_M03[1];
				11'd518:M <= line_M03[30];	11'd528:M <= line_M03[20];	11'd538:M <= line_M03[10];	11'd548:M <= line_M03[0];
				default:M <= 0;
			endcase
		11'd326:
			case (pixel_col)
				11'd509:M <= line_M04[39];	11'd519:M <= line_M04[29];	11'd529:M <= line_M04[19];	11'd539:M <= line_M04[9];
				11'd510:M <= line_M04[38];	11'd520:M <= line_M04[28];	11'd530:M <= line_M04[18];	11'd540:M <= line_M04[8];
				11'd511:M <= line_M04[37];	11'd521:M <= line_M04[27];	11'd531:M <= line_M04[17];	11'd541:M <= line_M04[7];
				11'd512:M <= line_M04[36];	11'd522:M <= line_M04[26];	11'd532:M <= line_M04[16];	11'd542:M <= line_M04[6];
				11'd513:M <= line_M04[35];	11'd523:M <= line_M04[25];	11'd533:M <= line_M04[15];	11'd543:M <= line_M04[5];
				11'd514:M <= line_M04[34];	11'd524:M <= line_M04[24];	11'd534:M <= line_M04[14];	11'd544:M <= line_M04[4];
				11'd515:M <= line_M04[33];	11'd525:M <= line_M04[23];	11'd535:M <= line_M04[13];	11'd545:M <= line_M04[3];
				11'd516:M <= line_M04[32];	11'd526:M <= line_M04[22];	11'd536:M <= line_M04[12];	11'd546:M <= line_M04[2];
				11'd517:M <= line_M04[31];	11'd527:M <= line_M04[21];	11'd537:M <= line_M04[11];	11'd547:M <= line_M04[1];
				11'd518:M <= line_M04[30];	11'd528:M <= line_M04[20];	11'd538:M <= line_M04[10];	11'd548:M <= line_M04[0];
				default:M <= 0;
			endcase
		11'd327:
			case (pixel_col)
				11'd509:M <= line_M05[39];	11'd519:M <= line_M05[29];	11'd529:M <= line_M05[19];	11'd539:M <= line_M05[9];
				11'd510:M <= line_M05[38];	11'd520:M <= line_M05[28];	11'd530:M <= line_M05[18];	11'd540:M <= line_M05[8];
				11'd511:M <= line_M05[37];	11'd521:M <= line_M05[27];	11'd531:M <= line_M05[17];	11'd541:M <= line_M05[7];
				11'd512:M <= line_M05[36];	11'd522:M <= line_M05[26];	11'd532:M <= line_M05[16];	11'd542:M <= line_M05[6];
				11'd513:M <= line_M05[35];	11'd523:M <= line_M05[25];	11'd533:M <= line_M05[15];	11'd543:M <= line_M05[5];
				11'd514:M <= line_M05[34];	11'd524:M <= line_M05[24];	11'd534:M <= line_M05[14];	11'd544:M <= line_M05[4];
				11'd515:M <= line_M05[33];	11'd525:M <= line_M05[23];	11'd535:M <= line_M05[13];	11'd545:M <= line_M05[3];
				11'd516:M <= line_M05[32];	11'd526:M <= line_M05[22];	11'd536:M <= line_M05[12];	11'd546:M <= line_M05[2];
				11'd517:M <= line_M05[31];	11'd527:M <= line_M05[21];	11'd537:M <= line_M05[11];	11'd547:M <= line_M05[1];
				11'd518:M <= line_M05[30];	11'd528:M <= line_M05[20];	11'd538:M <= line_M05[10];	11'd548:M <= line_M05[0];
				default:M <= 0;
			endcase
		11'd328:
			case (pixel_col)
				11'd509:M <= line_M06[39];	11'd519:M <= line_M06[29];	11'd529:M <= line_M06[19];	11'd539:M <= line_M06[9];
				11'd510:M <= line_M06[38];	11'd520:M <= line_M06[28];	11'd530:M <= line_M06[18];	11'd540:M <= line_M06[8];
				11'd511:M <= line_M06[37];	11'd521:M <= line_M06[27];	11'd531:M <= line_M06[17];	11'd541:M <= line_M06[7];
				11'd512:M <= line_M06[36];	11'd522:M <= line_M06[26];	11'd532:M <= line_M06[16];	11'd542:M <= line_M06[6];
				11'd513:M <= line_M06[35];	11'd523:M <= line_M06[25];	11'd533:M <= line_M06[15];	11'd543:M <= line_M06[5];
				11'd514:M <= line_M06[34];	11'd524:M <= line_M06[24];	11'd534:M <= line_M06[14];	11'd544:M <= line_M06[4];
				11'd515:M <= line_M06[33];	11'd525:M <= line_M06[23];	11'd535:M <= line_M06[13];	11'd545:M <= line_M06[3];
				11'd516:M <= line_M06[32];	11'd526:M <= line_M06[22];	11'd536:M <= line_M06[12];	11'd546:M <= line_M06[2];
				11'd517:M <= line_M06[31];	11'd527:M <= line_M06[21];	11'd537:M <= line_M06[11];	11'd547:M <= line_M06[1];
				11'd518:M <= line_M06[30];	11'd528:M <= line_M06[20];	11'd538:M <= line_M06[10];	11'd548:M <= line_M06[0];
				default:M <= 0;
			endcase
		11'd329:
			case (pixel_col)
				11'd509:M <= line_M07[39];	11'd519:M <= line_M07[29];	11'd529:M <= line_M07[19];	11'd539:M <= line_M07[9];
				11'd510:M <= line_M07[38];	11'd520:M <= line_M07[28];	11'd530:M <= line_M07[18];	11'd540:M <= line_M07[8];
				11'd511:M <= line_M07[37];	11'd521:M <= line_M07[27];	11'd531:M <= line_M07[17];	11'd541:M <= line_M07[7];
				11'd512:M <= line_M07[36];	11'd522:M <= line_M07[26];	11'd532:M <= line_M07[16];	11'd542:M <= line_M07[6];
				11'd513:M <= line_M07[35];	11'd523:M <= line_M07[25];	11'd533:M <= line_M07[15];	11'd543:M <= line_M07[5];
				11'd514:M <= line_M07[34];	11'd524:M <= line_M07[24];	11'd534:M <= line_M07[14];	11'd544:M <= line_M07[4];
				11'd515:M <= line_M07[33];	11'd525:M <= line_M07[23];	11'd535:M <= line_M07[13];	11'd545:M <= line_M07[3];
				11'd516:M <= line_M07[32];	11'd526:M <= line_M07[22];	11'd536:M <= line_M07[12];	11'd546:M <= line_M07[2];
				11'd517:M <= line_M07[31];	11'd527:M <= line_M07[21];	11'd537:M <= line_M07[11];	11'd547:M <= line_M07[1];
				11'd518:M <= line_M07[30];	11'd528:M <= line_M07[20];	11'd538:M <= line_M07[10];	11'd548:M <= line_M07[0];
				default:M <= 0;
			endcase
		11'd330:
			case (pixel_col)
				11'd509:M <= line_M08[39];	11'd519:M <= line_M08[29];	11'd529:M <= line_M08[19];	11'd539:M <= line_M08[9];
				11'd510:M <= line_M08[38];	11'd520:M <= line_M08[28];	11'd530:M <= line_M08[18];	11'd540:M <= line_M08[8];
				11'd511:M <= line_M08[37];	11'd521:M <= line_M08[27];	11'd531:M <= line_M08[17];	11'd541:M <= line_M08[7];
				11'd512:M <= line_M08[36];	11'd522:M <= line_M08[26];	11'd532:M <= line_M08[16];	11'd542:M <= line_M08[6];
				11'd513:M <= line_M08[35];	11'd523:M <= line_M08[25];	11'd533:M <= line_M08[15];	11'd543:M <= line_M08[5];
				11'd514:M <= line_M08[34];	11'd524:M <= line_M08[24];	11'd534:M <= line_M08[14];	11'd544:M <= line_M08[4];
				11'd515:M <= line_M08[33];	11'd525:M <= line_M08[23];	11'd535:M <= line_M08[13];	11'd545:M <= line_M08[3];
				11'd516:M <= line_M08[32];	11'd526:M <= line_M08[22];	11'd536:M <= line_M08[12];	11'd546:M <= line_M08[2];
				11'd517:M <= line_M08[31];	11'd527:M <= line_M08[21];	11'd537:M <= line_M08[11];	11'd547:M <= line_M08[1];
				11'd518:M <= line_M08[30];	11'd528:M <= line_M08[20];	11'd538:M <= line_M08[10];	11'd548:M <= line_M08[0];
				default:M <= 0;
			endcase
		11'd331:
			case (pixel_col)
				11'd509:M <= line_M09[39];	11'd519:M <= line_M09[29];	11'd529:M <= line_M09[19];	11'd539:M <= line_M09[9];
				11'd510:M <= line_M09[38];	11'd520:M <= line_M09[28];	11'd530:M <= line_M09[18];	11'd540:M <= line_M09[8];
				11'd511:M <= line_M09[37];	11'd521:M <= line_M09[27];	11'd531:M <= line_M09[17];	11'd541:M <= line_M09[7];
				11'd512:M <= line_M09[36];	11'd522:M <= line_M09[26];	11'd532:M <= line_M09[16];	11'd542:M <= line_M09[6];
				11'd513:M <= line_M09[35];	11'd523:M <= line_M09[25];	11'd533:M <= line_M09[15];	11'd543:M <= line_M09[5];
				11'd514:M <= line_M09[34];	11'd524:M <= line_M09[24];	11'd534:M <= line_M09[14];	11'd544:M <= line_M09[4];
				11'd515:M <= line_M09[33];	11'd525:M <= line_M09[23];	11'd535:M <= line_M09[13];	11'd545:M <= line_M09[3];
				11'd516:M <= line_M09[32];	11'd526:M <= line_M09[22];	11'd536:M <= line_M09[12];	11'd546:M <= line_M09[2];
				11'd517:M <= line_M09[31];	11'd527:M <= line_M09[21];	11'd537:M <= line_M09[11];	11'd547:M <= line_M09[1];
				11'd518:M <= line_M09[30];	11'd528:M <= line_M09[20];	11'd538:M <= line_M09[10];	11'd548:M <= line_M09[0];
				default:M <= 0;
			endcase
		11'd332:
			case (pixel_col)
				11'd509:M <= line_M10[39];	11'd519:M <= line_M10[29];	11'd529:M <= line_M10[19];	11'd539:M <= line_M10[9];
				11'd510:M <= line_M10[38];	11'd520:M <= line_M10[28];	11'd530:M <= line_M10[18];	11'd540:M <= line_M10[8];
				11'd511:M <= line_M10[37];	11'd521:M <= line_M10[27];	11'd531:M <= line_M10[17];	11'd541:M <= line_M10[7];
				11'd512:M <= line_M10[36];	11'd522:M <= line_M10[26];	11'd532:M <= line_M10[16];	11'd542:M <= line_M10[6];
				11'd513:M <= line_M10[35];	11'd523:M <= line_M10[25];	11'd533:M <= line_M10[15];	11'd543:M <= line_M10[5];
				11'd514:M <= line_M10[34];	11'd524:M <= line_M10[24];	11'd534:M <= line_M10[14];	11'd544:M <= line_M10[4];
				11'd515:M <= line_M10[33];	11'd525:M <= line_M10[23];	11'd535:M <= line_M10[13];	11'd545:M <= line_M10[3];
				11'd516:M <= line_M10[32];	11'd526:M <= line_M10[22];	11'd536:M <= line_M10[12];	11'd546:M <= line_M10[2];
				11'd517:M <= line_M10[31];	11'd527:M <= line_M10[21];	11'd537:M <= line_M10[11];	11'd547:M <= line_M10[1];
				11'd518:M <= line_M10[30];	11'd528:M <= line_M10[20];	11'd538:M <= line_M10[10];	11'd548:M <= line_M10[0];
				default:M <= 0;
			endcase
		11'd333:
			case (pixel_col)
				11'd509:M <= line_M11[39];	11'd519:M <= line_M11[29];	11'd529:M <= line_M11[19];	11'd539:M <= line_M11[9];
				11'd510:M <= line_M11[38];	11'd520:M <= line_M11[28];	11'd530:M <= line_M11[18];	11'd540:M <= line_M11[8];
				11'd511:M <= line_M11[37];	11'd521:M <= line_M11[27];	11'd531:M <= line_M11[17];	11'd541:M <= line_M11[7];
				11'd512:M <= line_M11[36];	11'd522:M <= line_M11[26];	11'd532:M <= line_M11[16];	11'd542:M <= line_M11[6];
				11'd513:M <= line_M11[35];	11'd523:M <= line_M11[25];	11'd533:M <= line_M11[15];	11'd543:M <= line_M11[5];
				11'd514:M <= line_M11[34];	11'd524:M <= line_M11[24];	11'd534:M <= line_M11[14];	11'd544:M <= line_M11[4];
				11'd515:M <= line_M11[33];	11'd525:M <= line_M11[23];	11'd535:M <= line_M11[13];	11'd545:M <= line_M11[3];
				11'd516:M <= line_M11[32];	11'd526:M <= line_M11[22];	11'd536:M <= line_M11[12];	11'd546:M <= line_M11[2];
				11'd517:M <= line_M11[31];	11'd527:M <= line_M11[21];	11'd537:M <= line_M11[11];	11'd547:M <= line_M11[1];
				11'd518:M <= line_M11[30];	11'd528:M <= line_M11[20];	11'd538:M <= line_M11[10];	11'd548:M <= line_M11[0];
				default:M <= 0;
			endcase
		11'd334:
			case (pixel_col)
				11'd509:M <= line_M12[39];	11'd519:M <= line_M12[29];	11'd529:M <= line_M12[19];	11'd539:M <= line_M12[9];
				11'd510:M <= line_M12[38];	11'd520:M <= line_M12[28];	11'd530:M <= line_M12[18];	11'd540:M <= line_M12[8];
				11'd511:M <= line_M12[37];	11'd521:M <= line_M12[27];	11'd531:M <= line_M12[17];	11'd541:M <= line_M12[7];
				11'd512:M <= line_M12[36];	11'd522:M <= line_M12[26];	11'd532:M <= line_M12[16];	11'd542:M <= line_M12[6];
				11'd513:M <= line_M12[35];	11'd523:M <= line_M12[25];	11'd533:M <= line_M12[15];	11'd543:M <= line_M12[5];
				11'd514:M <= line_M12[34];	11'd524:M <= line_M12[24];	11'd534:M <= line_M12[14];	11'd544:M <= line_M12[4];
				11'd515:M <= line_M12[33];	11'd525:M <= line_M12[23];	11'd535:M <= line_M12[13];	11'd545:M <= line_M12[3];
				11'd516:M <= line_M12[32];	11'd526:M <= line_M12[22];	11'd536:M <= line_M12[12];	11'd546:M <= line_M12[2];
				11'd517:M <= line_M12[31];	11'd527:M <= line_M12[21];	11'd537:M <= line_M12[11];	11'd547:M <= line_M12[1];
				11'd518:M <= line_M12[30];	11'd528:M <= line_M12[20];	11'd538:M <= line_M12[10];	11'd548:M <= line_M12[0];
				default:M <= 0;
			endcase
		11'd335:
			case (pixel_col)
				11'd509:M <= line_M13[39];	11'd519:M <= line_M13[29];	11'd529:M <= line_M13[19];	11'd539:M <= line_M13[9];
				11'd510:M <= line_M13[38];	11'd520:M <= line_M13[28];	11'd530:M <= line_M13[18];	11'd540:M <= line_M13[8];
				11'd511:M <= line_M13[37];	11'd521:M <= line_M13[27];	11'd531:M <= line_M13[17];	11'd541:M <= line_M13[7];
				11'd512:M <= line_M13[36];	11'd522:M <= line_M13[26];	11'd532:M <= line_M13[16];	11'd542:M <= line_M13[6];
				11'd513:M <= line_M13[35];	11'd523:M <= line_M13[25];	11'd533:M <= line_M13[15];	11'd543:M <= line_M13[5];
				11'd514:M <= line_M13[34];	11'd524:M <= line_M13[24];	11'd534:M <= line_M13[14];	11'd544:M <= line_M13[4];
				11'd515:M <= line_M13[33];	11'd525:M <= line_M13[23];	11'd535:M <= line_M13[13];	11'd545:M <= line_M13[3];
				11'd516:M <= line_M13[32];	11'd526:M <= line_M13[22];	11'd536:M <= line_M13[12];	11'd546:M <= line_M13[2];
				11'd517:M <= line_M13[31];	11'd527:M <= line_M13[21];	11'd537:M <= line_M13[11];	11'd547:M <= line_M13[1];
				11'd518:M <= line_M13[30];	11'd528:M <= line_M13[20];	11'd538:M <= line_M13[10];	11'd548:M <= line_M13[0];
				default:M <= 0;
			endcase
		11'd336:
			case (pixel_col)
				11'd509:M <= line_M14[39];	11'd519:M <= line_M14[29];	11'd529:M <= line_M14[19];	11'd539:M <= line_M14[9];
				11'd510:M <= line_M14[38];	11'd520:M <= line_M14[28];	11'd530:M <= line_M14[18];	11'd540:M <= line_M14[8];
				11'd511:M <= line_M14[37];	11'd521:M <= line_M14[27];	11'd531:M <= line_M14[17];	11'd541:M <= line_M14[7];
				11'd512:M <= line_M14[36];	11'd522:M <= line_M14[26];	11'd532:M <= line_M14[16];	11'd542:M <= line_M14[6];
				11'd513:M <= line_M14[35];	11'd523:M <= line_M14[25];	11'd533:M <= line_M14[15];	11'd543:M <= line_M14[5];
				11'd514:M <= line_M14[34];	11'd524:M <= line_M14[24];	11'd534:M <= line_M14[14];	11'd544:M <= line_M14[4];
				11'd515:M <= line_M14[33];	11'd525:M <= line_M14[23];	11'd535:M <= line_M14[13];	11'd545:M <= line_M14[3];
				11'd516:M <= line_M14[32];	11'd526:M <= line_M14[22];	11'd536:M <= line_M14[12];	11'd546:M <= line_M14[2];
				11'd517:M <= line_M14[31];	11'd527:M <= line_M14[21];	11'd537:M <= line_M14[11];	11'd547:M <= line_M14[1];
				11'd518:M <= line_M14[30];	11'd528:M <= line_M14[20];	11'd538:M <= line_M14[10];	11'd548:M <= line_M14[0];
				default:M <= 0;
			endcase
		11'd337:
			case (pixel_col)
				11'd509:M <= line_M15[39];	11'd519:M <= line_M15[29];	11'd529:M <= line_M15[19];	11'd539:M <= line_M15[9];
				11'd510:M <= line_M15[38];	11'd520:M <= line_M15[28];	11'd530:M <= line_M15[18];	11'd540:M <= line_M15[8];
				11'd511:M <= line_M15[37];	11'd521:M <= line_M15[27];	11'd531:M <= line_M15[17];	11'd541:M <= line_M15[7];
				11'd512:M <= line_M15[36];	11'd522:M <= line_M15[26];	11'd532:M <= line_M15[16];	11'd542:M <= line_M15[6];
				11'd513:M <= line_M15[35];	11'd523:M <= line_M15[25];	11'd533:M <= line_M15[15];	11'd543:M <= line_M15[5];
				11'd514:M <= line_M15[34];	11'd524:M <= line_M15[24];	11'd534:M <= line_M15[14];	11'd544:M <= line_M15[4];
				11'd515:M <= line_M15[33];	11'd525:M <= line_M15[23];	11'd535:M <= line_M15[13];	11'd545:M <= line_M15[3];
				11'd516:M <= line_M15[32];	11'd526:M <= line_M15[22];	11'd536:M <= line_M15[12];	11'd546:M <= line_M15[2];
				11'd517:M <= line_M15[31];	11'd527:M <= line_M15[21];	11'd537:M <= line_M15[11];	11'd547:M <= line_M15[1];
				11'd518:M <= line_M15[30];	11'd528:M <= line_M15[20];	11'd538:M <= line_M15[10];	11'd548:M <= line_M15[0];
				default:M <= 0;
			endcase
		default:M <= 0;
	endcase
end


always @(posedge clk) begin
	case (pixel_row)
		11'd323:
			case (pixel_col)
				11'd559:E <= line_E01[39];	11'd569:E <= line_E01[29];	11'd579:E <= line_E01[19];	11'd589:E <= line_E01[9];
				11'd560:E <= line_E01[38];	11'd570:E <= line_E01[28];	11'd580:E <= line_E01[18];	11'd590:E <= line_E01[8];
				11'd561:E <= line_E01[37];	11'd571:E <= line_E01[27];	11'd581:E <= line_E01[17];	11'd591:E <= line_E01[7];
				11'd562:E <= line_E01[36];	11'd572:E <= line_E01[26];	11'd582:E <= line_E01[16];	11'd592:E <= line_E01[6];
				11'd563:E <= line_E01[35];	11'd573:E <= line_E01[25];	11'd583:E <= line_E01[15];	11'd593:E <= line_E01[5];
				11'd564:E <= line_E01[34];	11'd574:E <= line_E01[24];	11'd584:E <= line_E01[14];	11'd594:E <= line_E01[4];
				11'd565:E <= line_E01[33];	11'd575:E <= line_E01[23];	11'd585:E <= line_E01[13];	11'd595:E <= line_E01[3];
				11'd566:E <= line_E01[32];	11'd576:E <= line_E01[22];	11'd586:E <= line_E01[12];	11'd596:E <= line_E01[2];
				11'd567:E <= line_E01[31];	11'd577:E <= line_E01[21];	11'd587:E <= line_E01[11];	11'd597:E <= line_E01[1];
				11'd568:E <= line_E01[30];	11'd578:E <= line_E01[20];	11'd588:E <= line_E01[10];	11'd598:E <= line_E01[0];
				default:E <= 0;
			endcase
		11'd324:
			case (pixel_col)
				11'd559:E <= line_E02[39];	11'd569:E <= line_E02[29];	11'd579:E <= line_E02[19];	11'd589:E <= line_E02[9];
				11'd560:E <= line_E02[38];	11'd570:E <= line_E02[28];	11'd580:E <= line_E02[18];	11'd590:E <= line_E02[8];
				11'd561:E <= line_E02[37];	11'd571:E <= line_E02[27];	11'd581:E <= line_E02[17];	11'd591:E <= line_E02[7];
				11'd562:E <= line_E02[36];	11'd572:E <= line_E02[26];	11'd582:E <= line_E02[16];	11'd592:E <= line_E02[6];
				11'd563:E <= line_E02[35];	11'd573:E <= line_E02[25];	11'd583:E <= line_E02[15];	11'd593:E <= line_E02[5];
				11'd564:E <= line_E02[34];	11'd574:E <= line_E02[24];	11'd584:E <= line_E02[14];	11'd594:E <= line_E02[4];
				11'd565:E <= line_E02[33];	11'd575:E <= line_E02[23];	11'd585:E <= line_E02[13];	11'd595:E <= line_E02[3];
				11'd566:E <= line_E02[32];	11'd576:E <= line_E02[22];	11'd586:E <= line_E02[12];	11'd596:E <= line_E02[2];
				11'd567:E <= line_E02[31];	11'd577:E <= line_E02[21];	11'd587:E <= line_E02[11];	11'd597:E <= line_E02[1];
				11'd568:E <= line_E02[30];	11'd578:E <= line_E02[20];	11'd588:E <= line_E02[10];	11'd598:E <= line_E02[0];
				default:E <= 0;
			endcase
		11'd325:
			case (pixel_col)
				11'd559:E <= line_E03[39];	11'd569:E <= line_E03[29];	11'd579:E <= line_E03[19];	11'd589:E <= line_E03[9];
				11'd560:E <= line_E03[38];	11'd570:E <= line_E03[28];	11'd580:E <= line_E03[18];	11'd590:E <= line_E03[8];
				11'd561:E <= line_E03[37];	11'd571:E <= line_E03[27];	11'd581:E <= line_E03[17];	11'd591:E <= line_E03[7];
				11'd562:E <= line_E03[36];	11'd572:E <= line_E03[26];	11'd582:E <= line_E03[16];	11'd592:E <= line_E03[6];
				11'd563:E <= line_E03[35];	11'd573:E <= line_E03[25];	11'd583:E <= line_E03[15];	11'd593:E <= line_E03[5];
				11'd564:E <= line_E03[34];	11'd574:E <= line_E03[24];	11'd584:E <= line_E03[14];	11'd594:E <= line_E03[4];
				11'd565:E <= line_E03[33];	11'd575:E <= line_E03[23];	11'd585:E <= line_E03[13];	11'd595:E <= line_E03[3];
				11'd566:E <= line_E03[32];	11'd576:E <= line_E03[22];	11'd586:E <= line_E03[12];	11'd596:E <= line_E03[2];
				11'd567:E <= line_E03[31];	11'd577:E <= line_E03[21];	11'd587:E <= line_E03[11];	11'd597:E <= line_E03[1];
				11'd568:E <= line_E03[30];	11'd578:E <= line_E03[20];	11'd588:E <= line_E03[10];	11'd598:E <= line_E03[0];
				default:E <= 0;
			endcase
		11'd326:
			case (pixel_col)
				11'd559:E <= line_E04[39];	11'd569:E <= line_E04[29];	11'd579:E <= line_E04[19];	11'd589:E <= line_E04[9];
				11'd560:E <= line_E04[38];	11'd570:E <= line_E04[28];	11'd580:E <= line_E04[18];	11'd590:E <= line_E04[8];
				11'd561:E <= line_E04[37];	11'd571:E <= line_E04[27];	11'd581:E <= line_E04[17];	11'd591:E <= line_E04[7];
				11'd562:E <= line_E04[36];	11'd572:E <= line_E04[26];	11'd582:E <= line_E04[16];	11'd592:E <= line_E04[6];
				11'd563:E <= line_E04[35];	11'd573:E <= line_E04[25];	11'd583:E <= line_E04[15];	11'd593:E <= line_E04[5];
				11'd564:E <= line_E04[34];	11'd574:E <= line_E04[24];	11'd584:E <= line_E04[14];	11'd594:E <= line_E04[4];
				11'd565:E <= line_E04[33];	11'd575:E <= line_E04[23];	11'd585:E <= line_E04[13];	11'd595:E <= line_E04[3];
				11'd566:E <= line_E04[32];	11'd576:E <= line_E04[22];	11'd586:E <= line_E04[12];	11'd596:E <= line_E04[2];
				11'd567:E <= line_E04[31];	11'd577:E <= line_E04[21];	11'd587:E <= line_E04[11];	11'd597:E <= line_E04[1];
				11'd568:E <= line_E04[30];	11'd578:E <= line_E04[20];	11'd588:E <= line_E04[10];	11'd598:E <= line_E04[0];
				default:E <= 0;
			endcase
		11'd327:
			case (pixel_col)
				11'd559:E <= line_E05[39];	11'd569:E <= line_E05[29];	11'd579:E <= line_E05[19];	11'd589:E <= line_E05[9];
				11'd560:E <= line_E05[38];	11'd570:E <= line_E05[28];	11'd580:E <= line_E05[18];	11'd590:E <= line_E05[8];
				11'd561:E <= line_E05[37];	11'd571:E <= line_E05[27];	11'd581:E <= line_E05[17];	11'd591:E <= line_E05[7];
				11'd562:E <= line_E05[36];	11'd572:E <= line_E05[26];	11'd582:E <= line_E05[16];	11'd592:E <= line_E05[6];
				11'd563:E <= line_E05[35];	11'd573:E <= line_E05[25];	11'd583:E <= line_E05[15];	11'd593:E <= line_E05[5];
				11'd564:E <= line_E05[34];	11'd574:E <= line_E05[24];	11'd584:E <= line_E05[14];	11'd594:E <= line_E05[4];
				11'd565:E <= line_E05[33];	11'd575:E <= line_E05[23];	11'd585:E <= line_E05[13];	11'd595:E <= line_E05[3];
				11'd566:E <= line_E05[32];	11'd576:E <= line_E05[22];	11'd586:E <= line_E05[12];	11'd596:E <= line_E05[2];
				11'd567:E <= line_E05[31];	11'd577:E <= line_E05[21];	11'd587:E <= line_E05[11];	11'd597:E <= line_E05[1];
				11'd568:E <= line_E05[30];	11'd578:E <= line_E05[20];	11'd588:E <= line_E05[10];	11'd598:E <= line_E05[0];
				default:E <= 0;
			endcase
		11'd328:
			case (pixel_col)
				11'd559:E <= line_E06[39];	11'd569:E <= line_E06[29];	11'd579:E <= line_E06[19];	11'd589:E <= line_E06[9];
				11'd560:E <= line_E06[38];	11'd570:E <= line_E06[28];	11'd580:E <= line_E06[18];	11'd590:E <= line_E06[8];
				11'd561:E <= line_E06[37];	11'd571:E <= line_E06[27];	11'd581:E <= line_E06[17];	11'd591:E <= line_E06[7];
				11'd562:E <= line_E06[36];	11'd572:E <= line_E06[26];	11'd582:E <= line_E06[16];	11'd592:E <= line_E06[6];
				11'd563:E <= line_E06[35];	11'd573:E <= line_E06[25];	11'd583:E <= line_E06[15];	11'd593:E <= line_E06[5];
				11'd564:E <= line_E06[34];	11'd574:E <= line_E06[24];	11'd584:E <= line_E06[14];	11'd594:E <= line_E06[4];
				11'd565:E <= line_E06[33];	11'd575:E <= line_E06[23];	11'd585:E <= line_E06[13];	11'd595:E <= line_E06[3];
				11'd566:E <= line_E06[32];	11'd576:E <= line_E06[22];	11'd586:E <= line_E06[12];	11'd596:E <= line_E06[2];
				11'd567:E <= line_E06[31];	11'd577:E <= line_E06[21];	11'd587:E <= line_E06[11];	11'd597:E <= line_E06[1];
				11'd568:E <= line_E06[30];	11'd578:E <= line_E06[20];	11'd588:E <= line_E06[10];	11'd598:E <= line_E06[0];
				default:E <= 0;
			endcase
		11'd329:
			case (pixel_col)
				11'd559:E <= line_E07[39];	11'd569:E <= line_E07[29];	11'd579:E <= line_E07[19];	11'd589:E <= line_E07[9];
				11'd560:E <= line_E07[38];	11'd570:E <= line_E07[28];	11'd580:E <= line_E07[18];	11'd590:E <= line_E07[8];
				11'd561:E <= line_E07[37];	11'd571:E <= line_E07[27];	11'd581:E <= line_E07[17];	11'd591:E <= line_E07[7];
				11'd562:E <= line_E07[36];	11'd572:E <= line_E07[26];	11'd582:E <= line_E07[16];	11'd592:E <= line_E07[6];
				11'd563:E <= line_E07[35];	11'd573:E <= line_E07[25];	11'd583:E <= line_E07[15];	11'd593:E <= line_E07[5];
				11'd564:E <= line_E07[34];	11'd574:E <= line_E07[24];	11'd584:E <= line_E07[14];	11'd594:E <= line_E07[4];
				11'd565:E <= line_E07[33];	11'd575:E <= line_E07[23];	11'd585:E <= line_E07[13];	11'd595:E <= line_E07[3];
				11'd566:E <= line_E07[32];	11'd576:E <= line_E07[22];	11'd586:E <= line_E07[12];	11'd596:E <= line_E07[2];
				11'd567:E <= line_E07[31];	11'd577:E <= line_E07[21];	11'd587:E <= line_E07[11];	11'd597:E <= line_E07[1];
				11'd568:E <= line_E07[30];	11'd578:E <= line_E07[20];	11'd588:E <= line_E07[10];	11'd598:E <= line_E07[0];
				default:E <= 0;
			endcase
		11'd330:
			case (pixel_col)
				11'd559:E <= line_E08[39];	11'd569:E <= line_E08[29];	11'd579:E <= line_E08[19];	11'd589:E <= line_E08[9];
				11'd560:E <= line_E08[38];	11'd570:E <= line_E08[28];	11'd580:E <= line_E08[18];	11'd590:E <= line_E08[8];
				11'd561:E <= line_E08[37];	11'd571:E <= line_E08[27];	11'd581:E <= line_E08[17];	11'd591:E <= line_E08[7];
				11'd562:E <= line_E08[36];	11'd572:E <= line_E08[26];	11'd582:E <= line_E08[16];	11'd592:E <= line_E08[6];
				11'd563:E <= line_E08[35];	11'd573:E <= line_E08[25];	11'd583:E <= line_E08[15];	11'd593:E <= line_E08[5];
				11'd564:E <= line_E08[34];	11'd574:E <= line_E08[24];	11'd584:E <= line_E08[14];	11'd594:E <= line_E08[4];
				11'd565:E <= line_E08[33];	11'd575:E <= line_E08[23];	11'd585:E <= line_E08[13];	11'd595:E <= line_E08[3];
				11'd566:E <= line_E08[32];	11'd576:E <= line_E08[22];	11'd586:E <= line_E08[12];	11'd596:E <= line_E08[2];
				11'd567:E <= line_E08[31];	11'd577:E <= line_E08[21];	11'd587:E <= line_E08[11];	11'd597:E <= line_E08[1];
				11'd568:E <= line_E08[30];	11'd578:E <= line_E08[20];	11'd588:E <= line_E08[10];	11'd598:E <= line_E08[0];
				default:E <= 0;
			endcase
		11'd331:
			case (pixel_col)
				11'd559:E <= line_E09[39];	11'd569:E <= line_E09[29];	11'd579:E <= line_E09[19];	11'd589:E <= line_E09[9];
				11'd560:E <= line_E09[38];	11'd570:E <= line_E09[28];	11'd580:E <= line_E09[18];	11'd590:E <= line_E09[8];
				11'd561:E <= line_E09[37];	11'd571:E <= line_E09[27];	11'd581:E <= line_E09[17];	11'd591:E <= line_E09[7];
				11'd562:E <= line_E09[36];	11'd572:E <= line_E09[26];	11'd582:E <= line_E09[16];	11'd592:E <= line_E09[6];
				11'd563:E <= line_E09[35];	11'd573:E <= line_E09[25];	11'd583:E <= line_E09[15];	11'd593:E <= line_E09[5];
				11'd564:E <= line_E09[34];	11'd574:E <= line_E09[24];	11'd584:E <= line_E09[14];	11'd594:E <= line_E09[4];
				11'd565:E <= line_E09[33];	11'd575:E <= line_E09[23];	11'd585:E <= line_E09[13];	11'd595:E <= line_E09[3];
				11'd566:E <= line_E09[32];	11'd576:E <= line_E09[22];	11'd586:E <= line_E09[12];	11'd596:E <= line_E09[2];
				11'd567:E <= line_E09[31];	11'd577:E <= line_E09[21];	11'd587:E <= line_E09[11];	11'd597:E <= line_E09[1];
				11'd568:E <= line_E09[30];	11'd578:E <= line_E09[20];	11'd588:E <= line_E09[10];	11'd598:E <= line_E09[0];
				default:E <= 0;
			endcase
		11'd332:
			case (pixel_col)
				11'd559:E <= line_E10[39];	11'd569:E <= line_E10[29];	11'd579:E <= line_E10[19];	11'd589:E <= line_E10[9];
				11'd560:E <= line_E10[38];	11'd570:E <= line_E10[28];	11'd580:E <= line_E10[18];	11'd590:E <= line_E10[8];
				11'd561:E <= line_E10[37];	11'd571:E <= line_E10[27];	11'd581:E <= line_E10[17];	11'd591:E <= line_E10[7];
				11'd562:E <= line_E10[36];	11'd572:E <= line_E10[26];	11'd582:E <= line_E10[16];	11'd592:E <= line_E10[6];
				11'd563:E <= line_E10[35];	11'd573:E <= line_E10[25];	11'd583:E <= line_E10[15];	11'd593:E <= line_E10[5];
				11'd564:E <= line_E10[34];	11'd574:E <= line_E10[24];	11'd584:E <= line_E10[14];	11'd594:E <= line_E10[4];
				11'd565:E <= line_E10[33];	11'd575:E <= line_E10[23];	11'd585:E <= line_E10[13];	11'd595:E <= line_E10[3];
				11'd566:E <= line_E10[32];	11'd576:E <= line_E10[22];	11'd586:E <= line_E10[12];	11'd596:E <= line_E10[2];
				11'd567:E <= line_E10[31];	11'd577:E <= line_E10[21];	11'd587:E <= line_E10[11];	11'd597:E <= line_E10[1];
				11'd568:E <= line_E10[30];	11'd578:E <= line_E10[20];	11'd588:E <= line_E10[10];	11'd598:E <= line_E10[0];
				default:E <= 0;
			endcase
		11'd333:
			case (pixel_col)
				11'd559:E <= line_E11[39];	11'd569:E <= line_E11[29];	11'd579:E <= line_E11[19];	11'd589:E <= line_E11[9];
				11'd560:E <= line_E11[38];	11'd570:E <= line_E11[28];	11'd580:E <= line_E11[18];	11'd590:E <= line_E11[8];
				11'd561:E <= line_E11[37];	11'd571:E <= line_E11[27];	11'd581:E <= line_E11[17];	11'd591:E <= line_E11[7];
				11'd562:E <= line_E11[36];	11'd572:E <= line_E11[26];	11'd582:E <= line_E11[16];	11'd592:E <= line_E11[6];
				11'd563:E <= line_E11[35];	11'd573:E <= line_E11[25];	11'd583:E <= line_E11[15];	11'd593:E <= line_E11[5];
				11'd564:E <= line_E11[34];	11'd574:E <= line_E11[24];	11'd584:E <= line_E11[14];	11'd594:E <= line_E11[4];
				11'd565:E <= line_E11[33];	11'd575:E <= line_E11[23];	11'd585:E <= line_E11[13];	11'd595:E <= line_E11[3];
				11'd566:E <= line_E11[32];	11'd576:E <= line_E11[22];	11'd586:E <= line_E11[12];	11'd596:E <= line_E11[2];
				11'd567:E <= line_E11[31];	11'd577:E <= line_E11[21];	11'd587:E <= line_E11[11];	11'd597:E <= line_E11[1];
				11'd568:E <= line_E11[30];	11'd578:E <= line_E11[20];	11'd588:E <= line_E11[10];	11'd598:E <= line_E11[0];
				default:E <= 0;
			endcase
		11'd334:
			case (pixel_col)
				11'd559:E <= line_E12[39];	11'd569:E <= line_E12[29];	11'd579:E <= line_E12[19];	11'd589:E <= line_E12[9];
				11'd560:E <= line_E12[38];	11'd570:E <= line_E12[28];	11'd580:E <= line_E12[18];	11'd590:E <= line_E12[8];
				11'd561:E <= line_E12[37];	11'd571:E <= line_E12[27];	11'd581:E <= line_E12[17];	11'd591:E <= line_E12[7];
				11'd562:E <= line_E12[36];	11'd572:E <= line_E12[26];	11'd582:E <= line_E12[16];	11'd592:E <= line_E12[6];
				11'd563:E <= line_E12[35];	11'd573:E <= line_E12[25];	11'd583:E <= line_E12[15];	11'd593:E <= line_E12[5];
				11'd564:E <= line_E12[34];	11'd574:E <= line_E12[24];	11'd584:E <= line_E12[14];	11'd594:E <= line_E12[4];
				11'd565:E <= line_E12[33];	11'd575:E <= line_E12[23];	11'd585:E <= line_E12[13];	11'd595:E <= line_E12[3];
				11'd566:E <= line_E12[32];	11'd576:E <= line_E12[22];	11'd586:E <= line_E12[12];	11'd596:E <= line_E12[2];
				11'd567:E <= line_E12[31];	11'd577:E <= line_E12[21];	11'd587:E <= line_E12[11];	11'd597:E <= line_E12[1];
				11'd568:E <= line_E12[30];	11'd578:E <= line_E12[20];	11'd588:E <= line_E12[10];	11'd598:E <= line_E12[0];
				default:E <= 0;
			endcase
		11'd335:
			case (pixel_col)
				11'd559:E <= line_E13[39];	11'd569:E <= line_E13[29];	11'd579:E <= line_E13[19];	11'd589:E <= line_E13[9];
				11'd560:E <= line_E13[38];	11'd570:E <= line_E13[28];	11'd580:E <= line_E13[18];	11'd590:E <= line_E13[8];
				11'd561:E <= line_E13[37];	11'd571:E <= line_E13[27];	11'd581:E <= line_E13[17];	11'd591:E <= line_E13[7];
				11'd562:E <= line_E13[36];	11'd572:E <= line_E13[26];	11'd582:E <= line_E13[16];	11'd592:E <= line_E13[6];
				11'd563:E <= line_E13[35];	11'd573:E <= line_E13[25];	11'd583:E <= line_E13[15];	11'd593:E <= line_E13[5];
				11'd564:E <= line_E13[34];	11'd574:E <= line_E13[24];	11'd584:E <= line_E13[14];	11'd594:E <= line_E13[4];
				11'd565:E <= line_E13[33];	11'd575:E <= line_E13[23];	11'd585:E <= line_E13[13];	11'd595:E <= line_E13[3];
				11'd566:E <= line_E13[32];	11'd576:E <= line_E13[22];	11'd586:E <= line_E13[12];	11'd596:E <= line_E13[2];
				11'd567:E <= line_E13[31];	11'd577:E <= line_E13[21];	11'd587:E <= line_E13[11];	11'd597:E <= line_E13[1];
				11'd568:E <= line_E13[30];	11'd578:E <= line_E13[20];	11'd588:E <= line_E13[10];	11'd598:E <= line_E13[0];
				default:E <= 0;
			endcase
		11'd336:
			case (pixel_col)
				11'd559:E <= line_E14[39];	11'd569:E <= line_E14[29];	11'd579:E <= line_E14[19];	11'd589:E <= line_E14[9];
				11'd560:E <= line_E14[38];	11'd570:E <= line_E14[28];	11'd580:E <= line_E14[18];	11'd590:E <= line_E14[8];
				11'd561:E <= line_E14[37];	11'd571:E <= line_E14[27];	11'd581:E <= line_E14[17];	11'd591:E <= line_E14[7];
				11'd562:E <= line_E14[36];	11'd572:E <= line_E14[26];	11'd582:E <= line_E14[16];	11'd592:E <= line_E14[6];
				11'd563:E <= line_E14[35];	11'd573:E <= line_E14[25];	11'd583:E <= line_E14[15];	11'd593:E <= line_E14[5];
				11'd564:E <= line_E14[34];	11'd574:E <= line_E14[24];	11'd584:E <= line_E14[14];	11'd594:E <= line_E14[4];
				11'd565:E <= line_E14[33];	11'd575:E <= line_E14[23];	11'd585:E <= line_E14[13];	11'd595:E <= line_E14[3];
				11'd566:E <= line_E14[32];	11'd576:E <= line_E14[22];	11'd586:E <= line_E14[12];	11'd596:E <= line_E14[2];
				11'd567:E <= line_E14[31];	11'd577:E <= line_E14[21];	11'd587:E <= line_E14[11];	11'd597:E <= line_E14[1];
				11'd568:E <= line_E14[30];	11'd578:E <= line_E14[20];	11'd588:E <= line_E14[10];	11'd598:E <= line_E14[0];
				default:E <= 0;
			endcase
		11'd337:
			case (pixel_col)
				11'd559:E <= line_E15[39];	11'd569:E <= line_E15[29];	11'd579:E <= line_E15[19];	11'd589:E <= line_E15[9];
				11'd560:E <= line_E15[38];	11'd570:E <= line_E15[28];	11'd580:E <= line_E15[18];	11'd590:E <= line_E15[8];
				11'd561:E <= line_E15[37];	11'd571:E <= line_E15[27];	11'd581:E <= line_E15[17];	11'd591:E <= line_E15[7];
				11'd562:E <= line_E15[36];	11'd572:E <= line_E15[26];	11'd582:E <= line_E15[16];	11'd592:E <= line_E15[6];
				11'd563:E <= line_E15[35];	11'd573:E <= line_E15[25];	11'd583:E <= line_E15[15];	11'd593:E <= line_E15[5];
				11'd564:E <= line_E15[34];	11'd574:E <= line_E15[24];	11'd584:E <= line_E15[14];	11'd594:E <= line_E15[4];
				11'd565:E <= line_E15[33];	11'd575:E <= line_E15[23];	11'd585:E <= line_E15[13];	11'd595:E <= line_E15[3];
				11'd566:E <= line_E15[32];	11'd576:E <= line_E15[22];	11'd586:E <= line_E15[12];	11'd596:E <= line_E15[2];
				11'd567:E <= line_E15[31];	11'd577:E <= line_E15[21];	11'd587:E <= line_E15[11];	11'd597:E <= line_E15[1];
				11'd568:E <= line_E15[30];	11'd578:E <= line_E15[20];	11'd588:E <= line_E15[10];	11'd598:E <= line_E15[0];
				default:E <= 0;
			endcase
		default:E <= 0;
	endcase
end

always @(posedge clk) begin
	case (pixel_row)
		11'd348:
			case (pixel_col)
				11'd409:O <= line_O01[39];	11'd419:O <= line_O01[29];	11'd429:O <= line_O01[19];	11'd439:O <= line_O01[9];
				11'd410:O <= line_O01[38];	11'd420:O <= line_O01[28];	11'd430:O <= line_O01[18];	11'd440:O <= line_O01[8];
				11'd411:O <= line_O01[37];	11'd421:O <= line_O01[27];	11'd431:O <= line_O01[17];	11'd441:O <= line_O01[7];
				11'd412:O <= line_O01[36];	11'd422:O <= line_O01[26];	11'd432:O <= line_O01[16];	11'd442:O <= line_O01[6];
				11'd413:O <= line_O01[35];	11'd423:O <= line_O01[25];	11'd433:O <= line_O01[15];	11'd443:O <= line_O01[5];
				11'd414:O <= line_O01[34];	11'd424:O <= line_O01[24];	11'd434:O <= line_O01[14];	11'd444:O <= line_O01[4];
				11'd415:O <= line_O01[33];	11'd425:O <= line_O01[23];	11'd435:O <= line_O01[13];	11'd445:O <= line_O01[3];
				11'd416:O <= line_O01[32];	11'd426:O <= line_O01[22];	11'd436:O <= line_O01[12];	11'd446:O <= line_O01[2];
				11'd417:O <= line_O01[31];	11'd427:O <= line_O01[21];	11'd437:O <= line_O01[11];	11'd447:O <= line_O01[1];
				11'd418:O <= line_O01[30];	11'd428:O <= line_O01[20];	11'd438:O <= line_O01[10];	11'd448:O <= line_O01[0];
				default:O <= 0;
			endcase
		11'd349:
			case (pixel_col)
				11'd409:O <= line_O02[39];	11'd419:O <= line_O02[29];	11'd429:O <= line_O02[19];	11'd439:O <= line_O02[9];
				11'd410:O <= line_O02[38];	11'd420:O <= line_O02[28];	11'd430:O <= line_O02[18];	11'd440:O <= line_O02[8];
				11'd411:O <= line_O02[37];	11'd421:O <= line_O02[27];	11'd431:O <= line_O02[17];	11'd441:O <= line_O02[7];
				11'd412:O <= line_O02[36];	11'd422:O <= line_O02[26];	11'd432:O <= line_O02[16];	11'd442:O <= line_O02[6];
				11'd413:O <= line_O02[35];	11'd423:O <= line_O02[25];	11'd433:O <= line_O02[15];	11'd443:O <= line_O02[5];
				11'd414:O <= line_O02[34];	11'd424:O <= line_O02[24];	11'd434:O <= line_O02[14];	11'd444:O <= line_O02[4];
				11'd415:O <= line_O02[33];	11'd425:O <= line_O02[23];	11'd435:O <= line_O02[13];	11'd445:O <= line_O02[3];
				11'd416:O <= line_O02[32];	11'd426:O <= line_O02[22];	11'd436:O <= line_O02[12];	11'd446:O <= line_O02[2];
				11'd417:O <= line_O02[31];	11'd427:O <= line_O02[21];	11'd437:O <= line_O02[11];	11'd447:O <= line_O02[1];
				11'd418:O <= line_O02[30];	11'd428:O <= line_O02[20];	11'd438:O <= line_O02[10];	11'd448:O <= line_O02[0];
				default:O <= 0;
			endcase
		11'd350:
			case (pixel_col)
				11'd409:O <= line_O03[39];	11'd419:O <= line_O03[29];	11'd429:O <= line_O03[19];	11'd439:O <= line_O03[9];
				11'd410:O <= line_O03[38];	11'd420:O <= line_O03[28];	11'd430:O <= line_O03[18];	11'd440:O <= line_O03[8];
				11'd411:O <= line_O03[37];	11'd421:O <= line_O03[27];	11'd431:O <= line_O03[17];	11'd441:O <= line_O03[7];
				11'd412:O <= line_O03[36];	11'd422:O <= line_O03[26];	11'd432:O <= line_O03[16];	11'd442:O <= line_O03[6];
				11'd413:O <= line_O03[35];	11'd423:O <= line_O03[25];	11'd433:O <= line_O03[15];	11'd443:O <= line_O03[5];
				11'd414:O <= line_O03[34];	11'd424:O <= line_O03[24];	11'd434:O <= line_O03[14];	11'd444:O <= line_O03[4];
				11'd415:O <= line_O03[33];	11'd425:O <= line_O03[23];	11'd435:O <= line_O03[13];	11'd445:O <= line_O03[3];
				11'd416:O <= line_O03[32];	11'd426:O <= line_O03[22];	11'd436:O <= line_O03[12];	11'd446:O <= line_O03[2];
				11'd417:O <= line_O03[31];	11'd427:O <= line_O03[21];	11'd437:O <= line_O03[11];	11'd447:O <= line_O03[1];
				11'd418:O <= line_O03[30];	11'd428:O <= line_O03[20];	11'd438:O <= line_O03[10];	11'd448:O <= line_O03[0];
				default:O <= 0;
			endcase
		11'd351:
			case (pixel_col)
				11'd409:O <= line_O04[39];	11'd419:O <= line_O04[29];	11'd429:O <= line_O04[19];	11'd439:O <= line_O04[9];
				11'd410:O <= line_O04[38];	11'd420:O <= line_O04[28];	11'd430:O <= line_O04[18];	11'd440:O <= line_O04[8];
				11'd411:O <= line_O04[37];	11'd421:O <= line_O04[27];	11'd431:O <= line_O04[17];	11'd441:O <= line_O04[7];
				11'd412:O <= line_O04[36];	11'd422:O <= line_O04[26];	11'd432:O <= line_O04[16];	11'd442:O <= line_O04[6];
				11'd413:O <= line_O04[35];	11'd423:O <= line_O04[25];	11'd433:O <= line_O04[15];	11'd443:O <= line_O04[5];
				11'd414:O <= line_O04[34];	11'd424:O <= line_O04[24];	11'd434:O <= line_O04[14];	11'd444:O <= line_O04[4];
				11'd415:O <= line_O04[33];	11'd425:O <= line_O04[23];	11'd435:O <= line_O04[13];	11'd445:O <= line_O04[3];
				11'd416:O <= line_O04[32];	11'd426:O <= line_O04[22];	11'd436:O <= line_O04[12];	11'd446:O <= line_O04[2];
				11'd417:O <= line_O04[31];	11'd427:O <= line_O04[21];	11'd437:O <= line_O04[11];	11'd447:O <= line_O04[1];
				11'd418:O <= line_O04[30];	11'd428:O <= line_O04[20];	11'd438:O <= line_O04[10];	11'd448:O <= line_O04[0];
				default:O <= 0;
			endcase
		11'd352:
			case (pixel_col)
				11'd409:O <= line_O05[39];	11'd419:O <= line_O05[29];	11'd429:O <= line_O05[19];	11'd439:O <= line_O05[9];
				11'd410:O <= line_O05[38];	11'd420:O <= line_O05[28];	11'd430:O <= line_O05[18];	11'd440:O <= line_O05[8];
				11'd411:O <= line_O05[37];	11'd421:O <= line_O05[27];	11'd431:O <= line_O05[17];	11'd441:O <= line_O05[7];
				11'd412:O <= line_O05[36];	11'd422:O <= line_O05[26];	11'd432:O <= line_O05[16];	11'd442:O <= line_O05[6];
				11'd413:O <= line_O05[35];	11'd423:O <= line_O05[25];	11'd433:O <= line_O05[15];	11'd443:O <= line_O05[5];
				11'd414:O <= line_O05[34];	11'd424:O <= line_O05[24];	11'd434:O <= line_O05[14];	11'd444:O <= line_O05[4];
				11'd415:O <= line_O05[33];	11'd425:O <= line_O05[23];	11'd435:O <= line_O05[13];	11'd445:O <= line_O05[3];
				11'd416:O <= line_O05[32];	11'd426:O <= line_O05[22];	11'd436:O <= line_O05[12];	11'd446:O <= line_O05[2];
				11'd417:O <= line_O05[31];	11'd427:O <= line_O05[21];	11'd437:O <= line_O05[11];	11'd447:O <= line_O05[1];
				11'd418:O <= line_O05[30];	11'd428:O <= line_O05[20];	11'd438:O <= line_O05[10];	11'd448:O <= line_O05[0];
				default:O <= 0;
			endcase
		11'd353:
			case (pixel_col)
				11'd409:O <= line_O06[39];	11'd419:O <= line_O06[29];	11'd429:O <= line_O06[19];	11'd439:O <= line_O06[9];
				11'd410:O <= line_O06[38];	11'd420:O <= line_O06[28];	11'd430:O <= line_O06[18];	11'd440:O <= line_O06[8];
				11'd411:O <= line_O06[37];	11'd421:O <= line_O06[27];	11'd431:O <= line_O06[17];	11'd441:O <= line_O06[7];
				11'd412:O <= line_O06[36];	11'd422:O <= line_O06[26];	11'd432:O <= line_O06[16];	11'd442:O <= line_O06[6];
				11'd413:O <= line_O06[35];	11'd423:O <= line_O06[25];	11'd433:O <= line_O06[15];	11'd443:O <= line_O06[5];
				11'd414:O <= line_O06[34];	11'd424:O <= line_O06[24];	11'd434:O <= line_O06[14];	11'd444:O <= line_O06[4];
				11'd415:O <= line_O06[33];	11'd425:O <= line_O06[23];	11'd435:O <= line_O06[13];	11'd445:O <= line_O06[3];
				11'd416:O <= line_O06[32];	11'd426:O <= line_O06[22];	11'd436:O <= line_O06[12];	11'd446:O <= line_O06[2];
				11'd417:O <= line_O06[31];	11'd427:O <= line_O06[21];	11'd437:O <= line_O06[11];	11'd447:O <= line_O06[1];
				11'd418:O <= line_O06[30];	11'd428:O <= line_O06[20];	11'd438:O <= line_O06[10];	11'd448:O <= line_O06[0];
				default:O <= 0;
			endcase
		11'd354:
			case (pixel_col)
				11'd409:O <= line_O07[39];	11'd419:O <= line_O07[29];	11'd429:O <= line_O07[19];	11'd439:O <= line_O07[9];
				11'd410:O <= line_O07[38];	11'd420:O <= line_O07[28];	11'd430:O <= line_O07[18];	11'd440:O <= line_O07[8];
				11'd411:O <= line_O07[37];	11'd421:O <= line_O07[27];	11'd431:O <= line_O07[17];	11'd441:O <= line_O07[7];
				11'd412:O <= line_O07[36];	11'd422:O <= line_O07[26];	11'd432:O <= line_O07[16];	11'd442:O <= line_O07[6];
				11'd413:O <= line_O07[35];	11'd423:O <= line_O07[25];	11'd433:O <= line_O07[15];	11'd443:O <= line_O07[5];
				11'd414:O <= line_O07[34];	11'd424:O <= line_O07[24];	11'd434:O <= line_O07[14];	11'd444:O <= line_O07[4];
				11'd415:O <= line_O07[33];	11'd425:O <= line_O07[23];	11'd435:O <= line_O07[13];	11'd445:O <= line_O07[3];
				11'd416:O <= line_O07[32];	11'd426:O <= line_O07[22];	11'd436:O <= line_O07[12];	11'd446:O <= line_O07[2];
				11'd417:O <= line_O07[31];	11'd427:O <= line_O07[21];	11'd437:O <= line_O07[11];	11'd447:O <= line_O07[1];
				11'd418:O <= line_O07[30];	11'd428:O <= line_O07[20];	11'd438:O <= line_O07[10];	11'd448:O <= line_O07[0];
				default:O <= 0;
			endcase
		11'd355:
			case (pixel_col)
				11'd409:O <= line_O08[39];	11'd419:O <= line_O08[29];	11'd429:O <= line_O08[19];	11'd439:O <= line_O08[9];
				11'd410:O <= line_O08[38];	11'd420:O <= line_O08[28];	11'd430:O <= line_O08[18];	11'd440:O <= line_O08[8];
				11'd411:O <= line_O08[37];	11'd421:O <= line_O08[27];	11'd431:O <= line_O08[17];	11'd441:O <= line_O08[7];
				11'd412:O <= line_O08[36];	11'd422:O <= line_O08[26];	11'd432:O <= line_O08[16];	11'd442:O <= line_O08[6];
				11'd413:O <= line_O08[35];	11'd423:O <= line_O08[25];	11'd433:O <= line_O08[15];	11'd443:O <= line_O08[5];
				11'd414:O <= line_O08[34];	11'd424:O <= line_O08[24];	11'd434:O <= line_O08[14];	11'd444:O <= line_O08[4];
				11'd415:O <= line_O08[33];	11'd425:O <= line_O08[23];	11'd435:O <= line_O08[13];	11'd445:O <= line_O08[3];
				11'd416:O <= line_O08[32];	11'd426:O <= line_O08[22];	11'd436:O <= line_O08[12];	11'd446:O <= line_O08[2];
				11'd417:O <= line_O08[31];	11'd427:O <= line_O08[21];	11'd437:O <= line_O08[11];	11'd447:O <= line_O08[1];
				11'd418:O <= line_O08[30];	11'd428:O <= line_O08[20];	11'd438:O <= line_O08[10];	11'd448:O <= line_O08[0];
				default:O <= 0;
			endcase
		11'd356:
			case (pixel_col)
				11'd409:O <= line_O09[39];	11'd419:O <= line_O09[29];	11'd429:O <= line_O09[19];	11'd439:O <= line_O09[9];
				11'd410:O <= line_O09[38];	11'd420:O <= line_O09[28];	11'd430:O <= line_O09[18];	11'd440:O <= line_O09[8];
				11'd411:O <= line_O09[37];	11'd421:O <= line_O09[27];	11'd431:O <= line_O09[17];	11'd441:O <= line_O09[7];
				11'd412:O <= line_O09[36];	11'd422:O <= line_O09[26];	11'd432:O <= line_O09[16];	11'd442:O <= line_O09[6];
				11'd413:O <= line_O09[35];	11'd423:O <= line_O09[25];	11'd433:O <= line_O09[15];	11'd443:O <= line_O09[5];
				11'd414:O <= line_O09[34];	11'd424:O <= line_O09[24];	11'd434:O <= line_O09[14];	11'd444:O <= line_O09[4];
				11'd415:O <= line_O09[33];	11'd425:O <= line_O09[23];	11'd435:O <= line_O09[13];	11'd445:O <= line_O09[3];
				11'd416:O <= line_O09[32];	11'd426:O <= line_O09[22];	11'd436:O <= line_O09[12];	11'd446:O <= line_O09[2];
				11'd417:O <= line_O09[31];	11'd427:O <= line_O09[21];	11'd437:O <= line_O09[11];	11'd447:O <= line_O09[1];
				11'd418:O <= line_O09[30];	11'd428:O <= line_O09[20];	11'd438:O <= line_O09[10];	11'd448:O <= line_O09[0];
				default:O <= 0;
			endcase
		11'd357:
			case (pixel_col)
				11'd409:O <= line_O10[39];	11'd419:O <= line_O10[29];	11'd429:O <= line_O10[19];	11'd439:O <= line_O10[9];
				11'd410:O <= line_O10[38];	11'd420:O <= line_O10[28];	11'd430:O <= line_O10[18];	11'd440:O <= line_O10[8];
				11'd411:O <= line_O10[37];	11'd421:O <= line_O10[27];	11'd431:O <= line_O10[17];	11'd441:O <= line_O10[7];
				11'd412:O <= line_O10[36];	11'd422:O <= line_O10[26];	11'd432:O <= line_O10[16];	11'd442:O <= line_O10[6];
				11'd413:O <= line_O10[35];	11'd423:O <= line_O10[25];	11'd433:O <= line_O10[15];	11'd443:O <= line_O10[5];
				11'd414:O <= line_O10[34];	11'd424:O <= line_O10[24];	11'd434:O <= line_O10[14];	11'd444:O <= line_O10[4];
				11'd415:O <= line_O10[33];	11'd425:O <= line_O10[23];	11'd435:O <= line_O10[13];	11'd445:O <= line_O10[3];
				11'd416:O <= line_O10[32];	11'd426:O <= line_O10[22];	11'd436:O <= line_O10[12];	11'd446:O <= line_O10[2];
				11'd417:O <= line_O10[31];	11'd427:O <= line_O10[21];	11'd437:O <= line_O10[11];	11'd447:O <= line_O10[1];
				11'd418:O <= line_O10[30];	11'd428:O <= line_O10[20];	11'd438:O <= line_O10[10];	11'd448:O <= line_O10[0];
				default:O <= 0;
			endcase
		11'd358:
			case (pixel_col)
				11'd409:O <= line_O11[39];	11'd419:O <= line_O11[29];	11'd429:O <= line_O11[19];	11'd439:O <= line_O11[9];
				11'd410:O <= line_O11[38];	11'd420:O <= line_O11[28];	11'd430:O <= line_O11[18];	11'd440:O <= line_O11[8];
				11'd411:O <= line_O11[37];	11'd421:O <= line_O11[27];	11'd431:O <= line_O11[17];	11'd441:O <= line_O11[7];
				11'd412:O <= line_O11[36];	11'd422:O <= line_O11[26];	11'd432:O <= line_O11[16];	11'd442:O <= line_O11[6];
				11'd413:O <= line_O11[35];	11'd423:O <= line_O11[25];	11'd433:O <= line_O11[15];	11'd443:O <= line_O11[5];
				11'd414:O <= line_O11[34];	11'd424:O <= line_O11[24];	11'd434:O <= line_O11[14];	11'd444:O <= line_O11[4];
				11'd415:O <= line_O11[33];	11'd425:O <= line_O11[23];	11'd435:O <= line_O11[13];	11'd445:O <= line_O11[3];
				11'd416:O <= line_O11[32];	11'd426:O <= line_O11[22];	11'd436:O <= line_O11[12];	11'd446:O <= line_O11[2];
				11'd417:O <= line_O11[31];	11'd427:O <= line_O11[21];	11'd437:O <= line_O11[11];	11'd447:O <= line_O11[1];
				11'd418:O <= line_O11[30];	11'd428:O <= line_O11[20];	11'd438:O <= line_O11[10];	11'd448:O <= line_O11[0];
				default:O <= 0;
			endcase
		11'd359:
			case (pixel_col)
				11'd409:O <= line_O12[39];	11'd419:O <= line_O12[29];	11'd429:O <= line_O12[19];	11'd439:O <= line_O12[9];
				11'd410:O <= line_O12[38];	11'd420:O <= line_O12[28];	11'd430:O <= line_O12[18];	11'd440:O <= line_O12[8];
				11'd411:O <= line_O12[37];	11'd421:O <= line_O12[27];	11'd431:O <= line_O12[17];	11'd441:O <= line_O12[7];
				11'd412:O <= line_O12[36];	11'd422:O <= line_O12[26];	11'd432:O <= line_O12[16];	11'd442:O <= line_O12[6];
				11'd413:O <= line_O12[35];	11'd423:O <= line_O12[25];	11'd433:O <= line_O12[15];	11'd443:O <= line_O12[5];
				11'd414:O <= line_O12[34];	11'd424:O <= line_O12[24];	11'd434:O <= line_O12[14];	11'd444:O <= line_O12[4];
				11'd415:O <= line_O12[33];	11'd425:O <= line_O12[23];	11'd435:O <= line_O12[13];	11'd445:O <= line_O12[3];
				11'd416:O <= line_O12[32];	11'd426:O <= line_O12[22];	11'd436:O <= line_O12[12];	11'd446:O <= line_O12[2];
				11'd417:O <= line_O12[31];	11'd427:O <= line_O12[21];	11'd437:O <= line_O12[11];	11'd447:O <= line_O12[1];
				11'd418:O <= line_O12[30];	11'd428:O <= line_O12[20];	11'd438:O <= line_O12[10];	11'd448:O <= line_O12[0];
				default:O <= 0;
			endcase
		11'd360:
			case (pixel_col)
				11'd409:O <= line_O13[39];	11'd419:O <= line_O13[29];	11'd429:O <= line_O13[19];	11'd439:O <= line_O13[9];
				11'd410:O <= line_O13[38];	11'd420:O <= line_O13[28];	11'd430:O <= line_O13[18];	11'd440:O <= line_O13[8];
				11'd411:O <= line_O13[37];	11'd421:O <= line_O13[27];	11'd431:O <= line_O13[17];	11'd441:O <= line_O13[7];
				11'd412:O <= line_O13[36];	11'd422:O <= line_O13[26];	11'd432:O <= line_O13[16];	11'd442:O <= line_O13[6];
				11'd413:O <= line_O13[35];	11'd423:O <= line_O13[25];	11'd433:O <= line_O13[15];	11'd443:O <= line_O13[5];
				11'd414:O <= line_O13[34];	11'd424:O <= line_O13[24];	11'd434:O <= line_O13[14];	11'd444:O <= line_O13[4];
				11'd415:O <= line_O13[33];	11'd425:O <= line_O13[23];	11'd435:O <= line_O13[13];	11'd445:O <= line_O13[3];
				11'd416:O <= line_O13[32];	11'd426:O <= line_O13[22];	11'd436:O <= line_O13[12];	11'd446:O <= line_O13[2];
				11'd417:O <= line_O13[31];	11'd427:O <= line_O13[21];	11'd437:O <= line_O13[11];	11'd447:O <= line_O13[1];
				11'd418:O <= line_O13[30];	11'd428:O <= line_O13[20];	11'd438:O <= line_O13[10];	11'd448:O <= line_O13[0];
				default:O <= 0;
			endcase
		11'd361:
			case (pixel_col)
				11'd409:O <= line_O14[39];	11'd419:O <= line_O14[29];	11'd429:O <= line_O14[19];	11'd439:O <= line_O14[9];
				11'd410:O <= line_O14[38];	11'd420:O <= line_O14[28];	11'd430:O <= line_O14[18];	11'd440:O <= line_O14[8];
				11'd411:O <= line_O14[37];	11'd421:O <= line_O14[27];	11'd431:O <= line_O14[17];	11'd441:O <= line_O14[7];
				11'd412:O <= line_O14[36];	11'd422:O <= line_O14[26];	11'd432:O <= line_O14[16];	11'd442:O <= line_O14[6];
				11'd413:O <= line_O14[35];	11'd423:O <= line_O14[25];	11'd433:O <= line_O14[15];	11'd443:O <= line_O14[5];
				11'd414:O <= line_O14[34];	11'd424:O <= line_O14[24];	11'd434:O <= line_O14[14];	11'd444:O <= line_O14[4];
				11'd415:O <= line_O14[33];	11'd425:O <= line_O14[23];	11'd435:O <= line_O14[13];	11'd445:O <= line_O14[3];
				11'd416:O <= line_O14[32];	11'd426:O <= line_O14[22];	11'd436:O <= line_O14[12];	11'd446:O <= line_O14[2];
				11'd417:O <= line_O14[31];	11'd427:O <= line_O14[21];	11'd437:O <= line_O14[11];	11'd447:O <= line_O14[1];
				11'd418:O <= line_O14[30];	11'd428:O <= line_O14[20];	11'd438:O <= line_O14[10];	11'd448:O <= line_O14[0];
				default:O <= 0;
			endcase
		11'd362:
			case (pixel_col)
				11'd409:O <= line_O15[39];	11'd419:O <= line_O15[29];	11'd429:O <= line_O15[19];	11'd439:O <= line_O15[9];
				11'd410:O <= line_O15[38];	11'd420:O <= line_O15[28];	11'd430:O <= line_O15[18];	11'd440:O <= line_O15[8];
				11'd411:O <= line_O15[37];	11'd421:O <= line_O15[27];	11'd431:O <= line_O15[17];	11'd441:O <= line_O15[7];
				11'd412:O <= line_O15[36];	11'd422:O <= line_O15[26];	11'd432:O <= line_O15[16];	11'd442:O <= line_O15[6];
				11'd413:O <= line_O15[35];	11'd423:O <= line_O15[25];	11'd433:O <= line_O15[15];	11'd443:O <= line_O15[5];
				11'd414:O <= line_O15[34];	11'd424:O <= line_O15[24];	11'd434:O <= line_O15[14];	11'd444:O <= line_O15[4];
				11'd415:O <= line_O15[33];	11'd425:O <= line_O15[23];	11'd435:O <= line_O15[13];	11'd445:O <= line_O15[3];
				11'd416:O <= line_O15[32];	11'd426:O <= line_O15[22];	11'd436:O <= line_O15[12];	11'd446:O <= line_O15[2];
				11'd417:O <= line_O15[31];	11'd427:O <= line_O15[21];	11'd437:O <= line_O15[11];	11'd447:O <= line_O15[1];
				11'd418:O <= line_O15[30];	11'd428:O <= line_O15[20];	11'd438:O <= line_O15[10];	11'd448:O <= line_O15[0];
				default:O <= 0;
			endcase
		default:O <= 0;
	endcase
end


always @(posedge clk) begin
	case (pixel_row)
		11'd348:
			case (pixel_col)
				11'd459:V <= line_V01[39];	11'd469:V <= line_V01[29];	11'd479:V <= line_V01[19];	11'd489:V <= line_V01[9];
				11'd460:V <= line_V01[38];	11'd470:V <= line_V01[28];	11'd480:V <= line_V01[18];	11'd490:V <= line_V01[8];
				11'd461:V <= line_V01[37];	11'd471:V <= line_V01[27];	11'd481:V <= line_V01[17];	11'd491:V <= line_V01[7];
				11'd462:V <= line_V01[36];	11'd472:V <= line_V01[26];	11'd482:V <= line_V01[16];	11'd492:V <= line_V01[6];
				11'd463:V <= line_V01[35];	11'd473:V <= line_V01[25];	11'd483:V <= line_V01[15];	11'd493:V <= line_V01[5];
				11'd464:V <= line_V01[34];	11'd474:V <= line_V01[24];	11'd484:V <= line_V01[14];	11'd494:V <= line_V01[4];
				11'd465:V <= line_V01[33];	11'd475:V <= line_V01[23];	11'd485:V <= line_V01[13];	11'd495:V <= line_V01[3];
				11'd466:V <= line_V01[32];	11'd476:V <= line_V01[22];	11'd486:V <= line_V01[12];	11'd496:V <= line_V01[2];
				11'd467:V <= line_V01[31];	11'd477:V <= line_V01[21];	11'd487:V <= line_V01[11];	11'd497:V <= line_V01[1];
				11'd468:V <= line_V01[30];	11'd478:V <= line_V01[20];	11'd488:V <= line_V01[10];	11'd498:V <= line_V01[0];
				default:V <= 0;
			endcase
		11'd349:
			case (pixel_col)
				11'd459:V <= line_V02[39];	11'd469:V <= line_V02[29];	11'd479:V <= line_V02[19];	11'd489:V <= line_V02[9];
				11'd460:V <= line_V02[38];	11'd470:V <= line_V02[28];	11'd480:V <= line_V02[18];	11'd490:V <= line_V02[8];
				11'd461:V <= line_V02[37];	11'd471:V <= line_V02[27];	11'd481:V <= line_V02[17];	11'd491:V <= line_V02[7];
				11'd462:V <= line_V02[36];	11'd472:V <= line_V02[26];	11'd482:V <= line_V02[16];	11'd492:V <= line_V02[6];
				11'd463:V <= line_V02[35];	11'd473:V <= line_V02[25];	11'd483:V <= line_V02[15];	11'd493:V <= line_V02[5];
				11'd464:V <= line_V02[34];	11'd474:V <= line_V02[24];	11'd484:V <= line_V02[14];	11'd494:V <= line_V02[4];
				11'd465:V <= line_V02[33];	11'd475:V <= line_V02[23];	11'd485:V <= line_V02[13];	11'd495:V <= line_V02[3];
				11'd466:V <= line_V02[32];	11'd476:V <= line_V02[22];	11'd486:V <= line_V02[12];	11'd496:V <= line_V02[2];
				11'd467:V <= line_V02[31];	11'd477:V <= line_V02[21];	11'd487:V <= line_V02[11];	11'd497:V <= line_V02[1];
				11'd468:V <= line_V02[30];	11'd478:V <= line_V02[20];	11'd488:V <= line_V02[10];	11'd498:V <= line_V02[0];
				default:V <= 0;
			endcase
		11'd350:
			case (pixel_col)
				11'd459:V <= line_V03[39];	11'd469:V <= line_V03[29];	11'd479:V <= line_V03[19];	11'd489:V <= line_V03[9];
				11'd460:V <= line_V03[38];	11'd470:V <= line_V03[28];	11'd480:V <= line_V03[18];	11'd490:V <= line_V03[8];
				11'd461:V <= line_V03[37];	11'd471:V <= line_V03[27];	11'd481:V <= line_V03[17];	11'd491:V <= line_V03[7];
				11'd462:V <= line_V03[36];	11'd472:V <= line_V03[26];	11'd482:V <= line_V03[16];	11'd492:V <= line_V03[6];
				11'd463:V <= line_V03[35];	11'd473:V <= line_V03[25];	11'd483:V <= line_V03[15];	11'd493:V <= line_V03[5];
				11'd464:V <= line_V03[34];	11'd474:V <= line_V03[24];	11'd484:V <= line_V03[14];	11'd494:V <= line_V03[4];
				11'd465:V <= line_V03[33];	11'd475:V <= line_V03[23];	11'd485:V <= line_V03[13];	11'd495:V <= line_V03[3];
				11'd466:V <= line_V03[32];	11'd476:V <= line_V03[22];	11'd486:V <= line_V03[12];	11'd496:V <= line_V03[2];
				11'd467:V <= line_V03[31];	11'd477:V <= line_V03[21];	11'd487:V <= line_V03[11];	11'd497:V <= line_V03[1];
				11'd468:V <= line_V03[30];	11'd478:V <= line_V03[20];	11'd488:V <= line_V03[10];	11'd498:V <= line_V03[0];
				default:V <= 0;
			endcase
		11'd351:
			case (pixel_col)
				11'd459:V <= line_V04[39];	11'd469:V <= line_V04[29];	11'd479:V <= line_V04[19];	11'd489:V <= line_V04[9];
				11'd460:V <= line_V04[38];	11'd470:V <= line_V04[28];	11'd480:V <= line_V04[18];	11'd490:V <= line_V04[8];
				11'd461:V <= line_V04[37];	11'd471:V <= line_V04[27];	11'd481:V <= line_V04[17];	11'd491:V <= line_V04[7];
				11'd462:V <= line_V04[36];	11'd472:V <= line_V04[26];	11'd482:V <= line_V04[16];	11'd492:V <= line_V04[6];
				11'd463:V <= line_V04[35];	11'd473:V <= line_V04[25];	11'd483:V <= line_V04[15];	11'd493:V <= line_V04[5];
				11'd464:V <= line_V04[34];	11'd474:V <= line_V04[24];	11'd484:V <= line_V04[14];	11'd494:V <= line_V04[4];
				11'd465:V <= line_V04[33];	11'd475:V <= line_V04[23];	11'd485:V <= line_V04[13];	11'd495:V <= line_V04[3];
				11'd466:V <= line_V04[32];	11'd476:V <= line_V04[22];	11'd486:V <= line_V04[12];	11'd496:V <= line_V04[2];
				11'd467:V <= line_V04[31];	11'd477:V <= line_V04[21];	11'd487:V <= line_V04[11];	11'd497:V <= line_V04[1];
				11'd468:V <= line_V04[30];	11'd478:V <= line_V04[20];	11'd488:V <= line_V04[10];	11'd498:V <= line_V04[0];
				default:V <= 0;
			endcase
		11'd352:
			case (pixel_col)
				11'd459:V <= line_V05[39];	11'd469:V <= line_V05[29];	11'd479:V <= line_V05[19];	11'd489:V <= line_V05[9];
				11'd460:V <= line_V05[38];	11'd470:V <= line_V05[28];	11'd480:V <= line_V05[18];	11'd490:V <= line_V05[8];
				11'd461:V <= line_V05[37];	11'd471:V <= line_V05[27];	11'd481:V <= line_V05[17];	11'd491:V <= line_V05[7];
				11'd462:V <= line_V05[36];	11'd472:V <= line_V05[26];	11'd482:V <= line_V05[16];	11'd492:V <= line_V05[6];
				11'd463:V <= line_V05[35];	11'd473:V <= line_V05[25];	11'd483:V <= line_V05[15];	11'd493:V <= line_V05[5];
				11'd464:V <= line_V05[34];	11'd474:V <= line_V05[24];	11'd484:V <= line_V05[14];	11'd494:V <= line_V05[4];
				11'd465:V <= line_V05[33];	11'd475:V <= line_V05[23];	11'd485:V <= line_V05[13];	11'd495:V <= line_V05[3];
				11'd466:V <= line_V05[32];	11'd476:V <= line_V05[22];	11'd486:V <= line_V05[12];	11'd496:V <= line_V05[2];
				11'd467:V <= line_V05[31];	11'd477:V <= line_V05[21];	11'd487:V <= line_V05[11];	11'd497:V <= line_V05[1];
				11'd468:V <= line_V05[30];	11'd478:V <= line_V05[20];	11'd488:V <= line_V05[10];	11'd498:V <= line_V05[0];
				default:V <= 0;
			endcase
		11'd353:
			case (pixel_col)
				11'd459:V <= line_V06[39];	11'd469:V <= line_V06[29];	11'd479:V <= line_V06[19];	11'd489:V <= line_V06[9];
				11'd460:V <= line_V06[38];	11'd470:V <= line_V06[28];	11'd480:V <= line_V06[18];	11'd490:V <= line_V06[8];
				11'd461:V <= line_V06[37];	11'd471:V <= line_V06[27];	11'd481:V <= line_V06[17];	11'd491:V <= line_V06[7];
				11'd462:V <= line_V06[36];	11'd472:V <= line_V06[26];	11'd482:V <= line_V06[16];	11'd492:V <= line_V06[6];
				11'd463:V <= line_V06[35];	11'd473:V <= line_V06[25];	11'd483:V <= line_V06[15];	11'd493:V <= line_V06[5];
				11'd464:V <= line_V06[34];	11'd474:V <= line_V06[24];	11'd484:V <= line_V06[14];	11'd494:V <= line_V06[4];
				11'd465:V <= line_V06[33];	11'd475:V <= line_V06[23];	11'd485:V <= line_V06[13];	11'd495:V <= line_V06[3];
				11'd466:V <= line_V06[32];	11'd476:V <= line_V06[22];	11'd486:V <= line_V06[12];	11'd496:V <= line_V06[2];
				11'd467:V <= line_V06[31];	11'd477:V <= line_V06[21];	11'd487:V <= line_V06[11];	11'd497:V <= line_V06[1];
				11'd468:V <= line_V06[30];	11'd478:V <= line_V06[20];	11'd488:V <= line_V06[10];	11'd498:V <= line_V06[0];
				default:V <= 0;
			endcase
		11'd354:
			case (pixel_col)
				11'd459:V <= line_V07[39];	11'd469:V <= line_V07[29];	11'd479:V <= line_V07[19];	11'd489:V <= line_V07[9];
				11'd460:V <= line_V07[38];	11'd470:V <= line_V07[28];	11'd480:V <= line_V07[18];	11'd490:V <= line_V07[8];
				11'd461:V <= line_V07[37];	11'd471:V <= line_V07[27];	11'd481:V <= line_V07[17];	11'd491:V <= line_V07[7];
				11'd462:V <= line_V07[36];	11'd472:V <= line_V07[26];	11'd482:V <= line_V07[16];	11'd492:V <= line_V07[6];
				11'd463:V <= line_V07[35];	11'd473:V <= line_V07[25];	11'd483:V <= line_V07[15];	11'd493:V <= line_V07[5];
				11'd464:V <= line_V07[34];	11'd474:V <= line_V07[24];	11'd484:V <= line_V07[14];	11'd494:V <= line_V07[4];
				11'd465:V <= line_V07[33];	11'd475:V <= line_V07[23];	11'd485:V <= line_V07[13];	11'd495:V <= line_V07[3];
				11'd466:V <= line_V07[32];	11'd476:V <= line_V07[22];	11'd486:V <= line_V07[12];	11'd496:V <= line_V07[2];
				11'd467:V <= line_V07[31];	11'd477:V <= line_V07[21];	11'd487:V <= line_V07[11];	11'd497:V <= line_V07[1];
				11'd468:V <= line_V07[30];	11'd478:V <= line_V07[20];	11'd488:V <= line_V07[10];	11'd498:V <= line_V07[0];
				default:V <= 0;
			endcase
		11'd355:
			case (pixel_col)
				11'd459:V <= line_V08[39];	11'd469:V <= line_V08[29];	11'd479:V <= line_V08[19];	11'd489:V <= line_V08[9];
				11'd460:V <= line_V08[38];	11'd470:V <= line_V08[28];	11'd480:V <= line_V08[18];	11'd490:V <= line_V08[8];
				11'd461:V <= line_V08[37];	11'd471:V <= line_V08[27];	11'd481:V <= line_V08[17];	11'd491:V <= line_V08[7];
				11'd462:V <= line_V08[36];	11'd472:V <= line_V08[26];	11'd482:V <= line_V08[16];	11'd492:V <= line_V08[6];
				11'd463:V <= line_V08[35];	11'd473:V <= line_V08[25];	11'd483:V <= line_V08[15];	11'd493:V <= line_V08[5];
				11'd464:V <= line_V08[34];	11'd474:V <= line_V08[24];	11'd484:V <= line_V08[14];	11'd494:V <= line_V08[4];
				11'd465:V <= line_V08[33];	11'd475:V <= line_V08[23];	11'd485:V <= line_V08[13];	11'd495:V <= line_V08[3];
				11'd466:V <= line_V08[32];	11'd476:V <= line_V08[22];	11'd486:V <= line_V08[12];	11'd496:V <= line_V08[2];
				11'd467:V <= line_V08[31];	11'd477:V <= line_V08[21];	11'd487:V <= line_V08[11];	11'd497:V <= line_V08[1];
				11'd468:V <= line_V08[30];	11'd478:V <= line_V08[20];	11'd488:V <= line_V08[10];	11'd498:V <= line_V08[0];
				default:V <= 0;
			endcase
		11'd356:
			case (pixel_col)
				11'd459:V <= line_V09[39];	11'd469:V <= line_V09[29];	11'd479:V <= line_V09[19];	11'd489:V <= line_V09[9];
				11'd460:V <= line_V09[38];	11'd470:V <= line_V09[28];	11'd480:V <= line_V09[18];	11'd490:V <= line_V09[8];
				11'd461:V <= line_V09[37];	11'd471:V <= line_V09[27];	11'd481:V <= line_V09[17];	11'd491:V <= line_V09[7];
				11'd462:V <= line_V09[36];	11'd472:V <= line_V09[26];	11'd482:V <= line_V09[16];	11'd492:V <= line_V09[6];
				11'd463:V <= line_V09[35];	11'd473:V <= line_V09[25];	11'd483:V <= line_V09[15];	11'd493:V <= line_V09[5];
				11'd464:V <= line_V09[34];	11'd474:V <= line_V09[24];	11'd484:V <= line_V09[14];	11'd494:V <= line_V09[4];
				11'd465:V <= line_V09[33];	11'd475:V <= line_V09[23];	11'd485:V <= line_V09[13];	11'd495:V <= line_V09[3];
				11'd466:V <= line_V09[32];	11'd476:V <= line_V09[22];	11'd486:V <= line_V09[12];	11'd496:V <= line_V09[2];
				11'd467:V <= line_V09[31];	11'd477:V <= line_V09[21];	11'd487:V <= line_V09[11];	11'd497:V <= line_V09[1];
				11'd468:V <= line_V09[30];	11'd478:V <= line_V09[20];	11'd488:V <= line_V09[10];	11'd498:V <= line_V09[0];
				default:V <= 0;
			endcase
		11'd357:
			case (pixel_col)
				11'd459:V <= line_V10[39];	11'd469:V <= line_V10[29];	11'd479:V <= line_V10[19];	11'd489:V <= line_V10[9];
				11'd460:V <= line_V10[38];	11'd470:V <= line_V10[28];	11'd480:V <= line_V10[18];	11'd490:V <= line_V10[8];
				11'd461:V <= line_V10[37];	11'd471:V <= line_V10[27];	11'd481:V <= line_V10[17];	11'd491:V <= line_V10[7];
				11'd462:V <= line_V10[36];	11'd472:V <= line_V10[26];	11'd482:V <= line_V10[16];	11'd492:V <= line_V10[6];
				11'd463:V <= line_V10[35];	11'd473:V <= line_V10[25];	11'd483:V <= line_V10[15];	11'd493:V <= line_V10[5];
				11'd464:V <= line_V10[34];	11'd474:V <= line_V10[24];	11'd484:V <= line_V10[14];	11'd494:V <= line_V10[4];
				11'd465:V <= line_V10[33];	11'd475:V <= line_V10[23];	11'd485:V <= line_V10[13];	11'd495:V <= line_V10[3];
				11'd466:V <= line_V10[32];	11'd476:V <= line_V10[22];	11'd486:V <= line_V10[12];	11'd496:V <= line_V10[2];
				11'd467:V <= line_V10[31];	11'd477:V <= line_V10[21];	11'd487:V <= line_V10[11];	11'd497:V <= line_V10[1];
				11'd468:V <= line_V10[30];	11'd478:V <= line_V10[20];	11'd488:V <= line_V10[10];	11'd498:V <= line_V10[0];
				default:V <= 0;
			endcase
		11'd358:
			case (pixel_col)
				11'd459:V <= line_V11[39];	11'd469:V <= line_V11[29];	11'd479:V <= line_V11[19];	11'd489:V <= line_V11[9];
				11'd460:V <= line_V11[38];	11'd470:V <= line_V11[28];	11'd480:V <= line_V11[18];	11'd490:V <= line_V11[8];
				11'd461:V <= line_V11[37];	11'd471:V <= line_V11[27];	11'd481:V <= line_V11[17];	11'd491:V <= line_V11[7];
				11'd462:V <= line_V11[36];	11'd472:V <= line_V11[26];	11'd482:V <= line_V11[16];	11'd492:V <= line_V11[6];
				11'd463:V <= line_V11[35];	11'd473:V <= line_V11[25];	11'd483:V <= line_V11[15];	11'd493:V <= line_V11[5];
				11'd464:V <= line_V11[34];	11'd474:V <= line_V11[24];	11'd484:V <= line_V11[14];	11'd494:V <= line_V11[4];
				11'd465:V <= line_V11[33];	11'd475:V <= line_V11[23];	11'd485:V <= line_V11[13];	11'd495:V <= line_V11[3];
				11'd466:V <= line_V11[32];	11'd476:V <= line_V11[22];	11'd486:V <= line_V11[12];	11'd496:V <= line_V11[2];
				11'd467:V <= line_V11[31];	11'd477:V <= line_V11[21];	11'd487:V <= line_V11[11];	11'd497:V <= line_V11[1];
				11'd468:V <= line_V11[30];	11'd478:V <= line_V11[20];	11'd488:V <= line_V11[10];	11'd498:V <= line_V11[0];
				default:V <= 0;
			endcase
		11'd359:
			case (pixel_col)
				11'd459:V <= line_V12[39];	11'd469:V <= line_V12[29];	11'd479:V <= line_V12[19];	11'd489:V <= line_V12[9];
				11'd460:V <= line_V12[38];	11'd470:V <= line_V12[28];	11'd480:V <= line_V12[18];	11'd490:V <= line_V12[8];
				11'd461:V <= line_V12[37];	11'd471:V <= line_V12[27];	11'd481:V <= line_V12[17];	11'd491:V <= line_V12[7];
				11'd462:V <= line_V12[36];	11'd472:V <= line_V12[26];	11'd482:V <= line_V12[16];	11'd492:V <= line_V12[6];
				11'd463:V <= line_V12[35];	11'd473:V <= line_V12[25];	11'd483:V <= line_V12[15];	11'd493:V <= line_V12[5];
				11'd464:V <= line_V12[34];	11'd474:V <= line_V12[24];	11'd484:V <= line_V12[14];	11'd494:V <= line_V12[4];
				11'd465:V <= line_V12[33];	11'd475:V <= line_V12[23];	11'd485:V <= line_V12[13];	11'd495:V <= line_V12[3];
				11'd466:V <= line_V12[32];	11'd476:V <= line_V12[22];	11'd486:V <= line_V12[12];	11'd496:V <= line_V12[2];
				11'd467:V <= line_V12[31];	11'd477:V <= line_V12[21];	11'd487:V <= line_V12[11];	11'd497:V <= line_V12[1];
				11'd468:V <= line_V12[30];	11'd478:V <= line_V12[20];	11'd488:V <= line_V12[10];	11'd498:V <= line_V12[0];
				default:V <= 0;
			endcase
		11'd360:
			case (pixel_col)
				11'd459:V <= line_V13[39];	11'd469:V <= line_V13[29];	11'd479:V <= line_V13[19];	11'd489:V <= line_V13[9];
				11'd460:V <= line_V13[38];	11'd470:V <= line_V13[28];	11'd480:V <= line_V13[18];	11'd490:V <= line_V13[8];
				11'd461:V <= line_V13[37];	11'd471:V <= line_V13[27];	11'd481:V <= line_V13[17];	11'd491:V <= line_V13[7];
				11'd462:V <= line_V13[36];	11'd472:V <= line_V13[26];	11'd482:V <= line_V13[16];	11'd492:V <= line_V13[6];
				11'd463:V <= line_V13[35];	11'd473:V <= line_V13[25];	11'd483:V <= line_V13[15];	11'd493:V <= line_V13[5];
				11'd464:V <= line_V13[34];	11'd474:V <= line_V13[24];	11'd484:V <= line_V13[14];	11'd494:V <= line_V13[4];
				11'd465:V <= line_V13[33];	11'd475:V <= line_V13[23];	11'd485:V <= line_V13[13];	11'd495:V <= line_V13[3];
				11'd466:V <= line_V13[32];	11'd476:V <= line_V13[22];	11'd486:V <= line_V13[12];	11'd496:V <= line_V13[2];
				11'd467:V <= line_V13[31];	11'd477:V <= line_V13[21];	11'd487:V <= line_V13[11];	11'd497:V <= line_V13[1];
				11'd468:V <= line_V13[30];	11'd478:V <= line_V13[20];	11'd488:V <= line_V13[10];	11'd498:V <= line_V13[0];
				default:V <= 0;
			endcase
		11'd361:
			case (pixel_col)
				11'd459:V <= line_V14[39];	11'd469:V <= line_V14[29];	11'd479:V <= line_V14[19];	11'd489:V <= line_V14[9];
				11'd460:V <= line_V14[38];	11'd470:V <= line_V14[28];	11'd480:V <= line_V14[18];	11'd490:V <= line_V14[8];
				11'd461:V <= line_V14[37];	11'd471:V <= line_V14[27];	11'd481:V <= line_V14[17];	11'd491:V <= line_V14[7];
				11'd462:V <= line_V14[36];	11'd472:V <= line_V14[26];	11'd482:V <= line_V14[16];	11'd492:V <= line_V14[6];
				11'd463:V <= line_V14[35];	11'd473:V <= line_V14[25];	11'd483:V <= line_V14[15];	11'd493:V <= line_V14[5];
				11'd464:V <= line_V14[34];	11'd474:V <= line_V14[24];	11'd484:V <= line_V14[14];	11'd494:V <= line_V14[4];
				11'd465:V <= line_V14[33];	11'd475:V <= line_V14[23];	11'd485:V <= line_V14[13];	11'd495:V <= line_V14[3];
				11'd466:V <= line_V14[32];	11'd476:V <= line_V14[22];	11'd486:V <= line_V14[12];	11'd496:V <= line_V14[2];
				11'd467:V <= line_V14[31];	11'd477:V <= line_V14[21];	11'd487:V <= line_V14[11];	11'd497:V <= line_V14[1];
				11'd468:V <= line_V14[30];	11'd478:V <= line_V14[20];	11'd488:V <= line_V14[10];	11'd498:V <= line_V14[0];
				default:V <= 0;
			endcase
		11'd362:
			case (pixel_col)
				11'd459:V <= line_V15[39];	11'd469:V <= line_V15[29];	11'd479:V <= line_V15[19];	11'd489:V <= line_V15[9];
				11'd460:V <= line_V15[38];	11'd470:V <= line_V15[28];	11'd480:V <= line_V15[18];	11'd490:V <= line_V15[8];
				11'd461:V <= line_V15[37];	11'd471:V <= line_V15[27];	11'd481:V <= line_V15[17];	11'd491:V <= line_V15[7];
				11'd462:V <= line_V15[36];	11'd472:V <= line_V15[26];	11'd482:V <= line_V15[16];	11'd492:V <= line_V15[6];
				11'd463:V <= line_V15[35];	11'd473:V <= line_V15[25];	11'd483:V <= line_V15[15];	11'd493:V <= line_V15[5];
				11'd464:V <= line_V15[34];	11'd474:V <= line_V15[24];	11'd484:V <= line_V15[14];	11'd494:V <= line_V15[4];
				11'd465:V <= line_V15[33];	11'd475:V <= line_V15[23];	11'd485:V <= line_V15[13];	11'd495:V <= line_V15[3];
				11'd466:V <= line_V15[32];	11'd476:V <= line_V15[22];	11'd486:V <= line_V15[12];	11'd496:V <= line_V15[2];
				11'd467:V <= line_V15[31];	11'd477:V <= line_V15[21];	11'd487:V <= line_V15[11];	11'd497:V <= line_V15[1];
				11'd468:V <= line_V15[30];	11'd478:V <= line_V15[20];	11'd488:V <= line_V15[10];	11'd498:V <= line_V15[0];
				default:V <= 0;
			endcase
		default:V <= 0;
	endcase
end


always @(posedge clk) begin
	case (pixel_row)
		11'd348:
			case (pixel_col)
				11'd509:E2 <= line_E01[39];	11'd519:E2 <= line_E01[29];	11'd529:E2 <= line_E01[19];	11'd539:E2 <= line_E01[9];
				11'd510:E2 <= line_E01[38];	11'd520:E2 <= line_E01[28];	11'd530:E2 <= line_E01[18];	11'd540:E2 <= line_E01[8];
				11'd511:E2 <= line_E01[37];	11'd521:E2 <= line_E01[27];	11'd531:E2 <= line_E01[17];	11'd541:E2 <= line_E01[7];
				11'd512:E2 <= line_E01[36];	11'd522:E2 <= line_E01[26];	11'd532:E2 <= line_E01[16];	11'd542:E2 <= line_E01[6];
				11'd513:E2 <= line_E01[35];	11'd523:E2 <= line_E01[25];	11'd533:E2 <= line_E01[15];	11'd543:E2 <= line_E01[5];
				11'd514:E2 <= line_E01[34];	11'd524:E2 <= line_E01[24];	11'd534:E2 <= line_E01[14];	11'd544:E2 <= line_E01[4];
				11'd515:E2 <= line_E01[33];	11'd525:E2 <= line_E01[23];	11'd535:E2 <= line_E01[13];	11'd545:E2 <= line_E01[3];
				11'd516:E2 <= line_E01[32];	11'd526:E2 <= line_E01[22];	11'd536:E2 <= line_E01[12];	11'd546:E2 <= line_E01[2];
				11'd517:E2 <= line_E01[31];	11'd527:E2 <= line_E01[21];	11'd537:E2 <= line_E01[11];	11'd547:E2 <= line_E01[1];
				11'd518:E2 <= line_E01[30];	11'd528:E2 <= line_E01[20];	11'd538:E2 <= line_E01[10];	11'd548:E2 <= line_E01[0];
				default:E2 <= 0;
			endcase
		11'd349:
			case (pixel_col)
				11'd509:E2 <= line_E02[39];	11'd519:E2 <= line_E02[29];	11'd529:E2 <= line_E02[19];	11'd539:E2 <= line_E02[9];
				11'd510:E2 <= line_E02[38];	11'd520:E2 <= line_E02[28];	11'd530:E2 <= line_E02[18];	11'd540:E2 <= line_E02[8];
				11'd511:E2 <= line_E02[37];	11'd521:E2 <= line_E02[27];	11'd531:E2 <= line_E02[17];	11'd541:E2 <= line_E02[7];
				11'd512:E2 <= line_E02[36];	11'd522:E2 <= line_E02[26];	11'd532:E2 <= line_E02[16];	11'd542:E2 <= line_E02[6];
				11'd513:E2 <= line_E02[35];	11'd523:E2 <= line_E02[25];	11'd533:E2 <= line_E02[15];	11'd543:E2 <= line_E02[5];
				11'd514:E2 <= line_E02[34];	11'd524:E2 <= line_E02[24];	11'd534:E2 <= line_E02[14];	11'd544:E2 <= line_E02[4];
				11'd515:E2 <= line_E02[33];	11'd525:E2 <= line_E02[23];	11'd535:E2 <= line_E02[13];	11'd545:E2 <= line_E02[3];
				11'd516:E2 <= line_E02[32];	11'd526:E2 <= line_E02[22];	11'd536:E2 <= line_E02[12];	11'd546:E2 <= line_E02[2];
				11'd517:E2 <= line_E02[31];	11'd527:E2 <= line_E02[21];	11'd537:E2 <= line_E02[11];	11'd547:E2 <= line_E02[1];
				11'd518:E2 <= line_E02[30];	11'd528:E2 <= line_E02[20];	11'd538:E2 <= line_E02[10];	11'd548:E2 <= line_E02[0];
				default:E2 <= 0;
			endcase
		11'd350:
			case (pixel_col)
				11'd509:E2 <= line_E03[39];	11'd519:E2 <= line_E03[29];	11'd529:E2 <= line_E03[19];	11'd539:E2 <= line_E03[9];
				11'd510:E2 <= line_E03[38];	11'd520:E2 <= line_E03[28];	11'd530:E2 <= line_E03[18];	11'd540:E2 <= line_E03[8];
				11'd511:E2 <= line_E03[37];	11'd521:E2 <= line_E03[27];	11'd531:E2 <= line_E03[17];	11'd541:E2 <= line_E03[7];
				11'd512:E2 <= line_E03[36];	11'd522:E2 <= line_E03[26];	11'd532:E2 <= line_E03[16];	11'd542:E2 <= line_E03[6];
				11'd513:E2 <= line_E03[35];	11'd523:E2 <= line_E03[25];	11'd533:E2 <= line_E03[15];	11'd543:E2 <= line_E03[5];
				11'd514:E2 <= line_E03[34];	11'd524:E2 <= line_E03[24];	11'd534:E2 <= line_E03[14];	11'd544:E2 <= line_E03[4];
				11'd515:E2 <= line_E03[33];	11'd525:E2 <= line_E03[23];	11'd535:E2 <= line_E03[13];	11'd545:E2 <= line_E03[3];
				11'd516:E2 <= line_E03[32];	11'd526:E2 <= line_E03[22];	11'd536:E2 <= line_E03[12];	11'd546:E2 <= line_E03[2];
				11'd517:E2 <= line_E03[31];	11'd527:E2 <= line_E03[21];	11'd537:E2 <= line_E03[11];	11'd547:E2 <= line_E03[1];
				11'd518:E2 <= line_E03[30];	11'd528:E2 <= line_E03[20];	11'd538:E2 <= line_E03[10];	11'd548:E2 <= line_E03[0];
				default:E2 <= 0;
			endcase
		11'd351:
			case (pixel_col)
				11'd509:E2 <= line_E04[39];	11'd519:E2 <= line_E04[29];	11'd529:E2 <= line_E04[19];	11'd539:E2 <= line_E04[9];
				11'd510:E2 <= line_E04[38];	11'd520:E2 <= line_E04[28];	11'd530:E2 <= line_E04[18];	11'd540:E2 <= line_E04[8];
				11'd511:E2 <= line_E04[37];	11'd521:E2 <= line_E04[27];	11'd531:E2 <= line_E04[17];	11'd541:E2 <= line_E04[7];
				11'd512:E2 <= line_E04[36];	11'd522:E2 <= line_E04[26];	11'd532:E2 <= line_E04[16];	11'd542:E2 <= line_E04[6];
				11'd513:E2 <= line_E04[35];	11'd523:E2 <= line_E04[25];	11'd533:E2 <= line_E04[15];	11'd543:E2 <= line_E04[5];
				11'd514:E2 <= line_E04[34];	11'd524:E2 <= line_E04[24];	11'd534:E2 <= line_E04[14];	11'd544:E2 <= line_E04[4];
				11'd515:E2 <= line_E04[33];	11'd525:E2 <= line_E04[23];	11'd535:E2 <= line_E04[13];	11'd545:E2 <= line_E04[3];
				11'd516:E2 <= line_E04[32];	11'd526:E2 <= line_E04[22];	11'd536:E2 <= line_E04[12];	11'd546:E2 <= line_E04[2];
				11'd517:E2 <= line_E04[31];	11'd527:E2 <= line_E04[21];	11'd537:E2 <= line_E04[11];	11'd547:E2 <= line_E04[1];
				11'd518:E2 <= line_E04[30];	11'd528:E2 <= line_E04[20];	11'd538:E2 <= line_E04[10];	11'd548:E2 <= line_E04[0];
				default:E2 <= 0;
			endcase
		11'd352:
			case (pixel_col)
				11'd509:E2 <= line_E05[39];	11'd519:E2 <= line_E05[29];	11'd529:E2 <= line_E05[19];	11'd539:E2 <= line_E05[9];
				11'd510:E2 <= line_E05[38];	11'd520:E2 <= line_E05[28];	11'd530:E2 <= line_E05[18];	11'd540:E2 <= line_E05[8];
				11'd511:E2 <= line_E05[37];	11'd521:E2 <= line_E05[27];	11'd531:E2 <= line_E05[17];	11'd541:E2 <= line_E05[7];
				11'd512:E2 <= line_E05[36];	11'd522:E2 <= line_E05[26];	11'd532:E2 <= line_E05[16];	11'd542:E2 <= line_E05[6];
				11'd513:E2 <= line_E05[35];	11'd523:E2 <= line_E05[25];	11'd533:E2 <= line_E05[15];	11'd543:E2 <= line_E05[5];
				11'd514:E2 <= line_E05[34];	11'd524:E2 <= line_E05[24];	11'd534:E2 <= line_E05[14];	11'd544:E2 <= line_E05[4];
				11'd515:E2 <= line_E05[33];	11'd525:E2 <= line_E05[23];	11'd535:E2 <= line_E05[13];	11'd545:E2 <= line_E05[3];
				11'd516:E2 <= line_E05[32];	11'd526:E2 <= line_E05[22];	11'd536:E2 <= line_E05[12];	11'd546:E2 <= line_E05[2];
				11'd517:E2 <= line_E05[31];	11'd527:E2 <= line_E05[21];	11'd537:E2 <= line_E05[11];	11'd547:E2 <= line_E05[1];
				11'd518:E2 <= line_E05[30];	11'd528:E2 <= line_E05[20];	11'd538:E2 <= line_E05[10];	11'd548:E2 <= line_E05[0];
				default:E2 <= 0;
			endcase
		11'd353:
			case (pixel_col)
				11'd509:E2 <= line_E06[39];	11'd519:E2 <= line_E06[29];	11'd529:E2 <= line_E06[19];	11'd539:E2 <= line_E06[9];
				11'd510:E2 <= line_E06[38];	11'd520:E2 <= line_E06[28];	11'd530:E2 <= line_E06[18];	11'd540:E2 <= line_E06[8];
				11'd511:E2 <= line_E06[37];	11'd521:E2 <= line_E06[27];	11'd531:E2 <= line_E06[17];	11'd541:E2 <= line_E06[7];
				11'd512:E2 <= line_E06[36];	11'd522:E2 <= line_E06[26];	11'd532:E2 <= line_E06[16];	11'd542:E2 <= line_E06[6];
				11'd513:E2 <= line_E06[35];	11'd523:E2 <= line_E06[25];	11'd533:E2 <= line_E06[15];	11'd543:E2 <= line_E06[5];
				11'd514:E2 <= line_E06[34];	11'd524:E2 <= line_E06[24];	11'd534:E2 <= line_E06[14];	11'd544:E2 <= line_E06[4];
				11'd515:E2 <= line_E06[33];	11'd525:E2 <= line_E06[23];	11'd535:E2 <= line_E06[13];	11'd545:E2 <= line_E06[3];
				11'd516:E2 <= line_E06[32];	11'd526:E2 <= line_E06[22];	11'd536:E2 <= line_E06[12];	11'd546:E2 <= line_E06[2];
				11'd517:E2 <= line_E06[31];	11'd527:E2 <= line_E06[21];	11'd537:E2 <= line_E06[11];	11'd547:E2 <= line_E06[1];
				11'd518:E2 <= line_E06[30];	11'd528:E2 <= line_E06[20];	11'd538:E2 <= line_E06[10];	11'd548:E2 <= line_E06[0];
				default:E2 <= 0;
			endcase
		11'd354:
			case (pixel_col)
				11'd509:E2 <= line_E07[39];	11'd519:E2 <= line_E07[29];	11'd529:E2 <= line_E07[19];	11'd539:E2 <= line_E07[9];
				11'd510:E2 <= line_E07[38];	11'd520:E2 <= line_E07[28];	11'd530:E2 <= line_E07[18];	11'd540:E2 <= line_E07[8];
				11'd511:E2 <= line_E07[37];	11'd521:E2 <= line_E07[27];	11'd531:E2 <= line_E07[17];	11'd541:E2 <= line_E07[7];
				11'd512:E2 <= line_E07[36];	11'd522:E2 <= line_E07[26];	11'd532:E2 <= line_E07[16];	11'd542:E2 <= line_E07[6];
				11'd513:E2 <= line_E07[35];	11'd523:E2 <= line_E07[25];	11'd533:E2 <= line_E07[15];	11'd543:E2 <= line_E07[5];
				11'd514:E2 <= line_E07[34];	11'd524:E2 <= line_E07[24];	11'd534:E2 <= line_E07[14];	11'd544:E2 <= line_E07[4];
				11'd515:E2 <= line_E07[33];	11'd525:E2 <= line_E07[23];	11'd535:E2 <= line_E07[13];	11'd545:E2 <= line_E07[3];
				11'd516:E2 <= line_E07[32];	11'd526:E2 <= line_E07[22];	11'd536:E2 <= line_E07[12];	11'd546:E2 <= line_E07[2];
				11'd517:E2 <= line_E07[31];	11'd527:E2 <= line_E07[21];	11'd537:E2 <= line_E07[11];	11'd547:E2 <= line_E07[1];
				11'd518:E2 <= line_E07[30];	11'd528:E2 <= line_E07[20];	11'd538:E2 <= line_E07[10];	11'd548:E2 <= line_E07[0];
				default:E2 <= 0;
			endcase
		11'd355:
			case (pixel_col)
				11'd509:E2 <= line_E08[39];	11'd519:E2 <= line_E08[29];	11'd529:E2 <= line_E08[19];	11'd539:E2 <= line_E08[9];
				11'd510:E2 <= line_E08[38];	11'd520:E2 <= line_E08[28];	11'd530:E2 <= line_E08[18];	11'd540:E2 <= line_E08[8];
				11'd511:E2 <= line_E08[37];	11'd521:E2 <= line_E08[27];	11'd531:E2 <= line_E08[17];	11'd541:E2 <= line_E08[7];
				11'd512:E2 <= line_E08[36];	11'd522:E2 <= line_E08[26];	11'd532:E2 <= line_E08[16];	11'd542:E2 <= line_E08[6];
				11'd513:E2 <= line_E08[35];	11'd523:E2 <= line_E08[25];	11'd533:E2 <= line_E08[15];	11'd543:E2 <= line_E08[5];
				11'd514:E2 <= line_E08[34];	11'd524:E2 <= line_E08[24];	11'd534:E2 <= line_E08[14];	11'd544:E2 <= line_E08[4];
				11'd515:E2 <= line_E08[33];	11'd525:E2 <= line_E08[23];	11'd535:E2 <= line_E08[13];	11'd545:E2 <= line_E08[3];
				11'd516:E2 <= line_E08[32];	11'd526:E2 <= line_E08[22];	11'd536:E2 <= line_E08[12];	11'd546:E2 <= line_E08[2];
				11'd517:E2 <= line_E08[31];	11'd527:E2 <= line_E08[21];	11'd537:E2 <= line_E08[11];	11'd547:E2 <= line_E08[1];
				11'd518:E2 <= line_E08[30];	11'd528:E2 <= line_E08[20];	11'd538:E2 <= line_E08[10];	11'd548:E2 <= line_E08[0];
				default:E2 <= 0;
			endcase
		11'd356:
			case (pixel_col)
				11'd509:E2 <= line_E09[39];	11'd519:E2 <= line_E09[29];	11'd529:E2 <= line_E09[19];	11'd539:E2 <= line_E09[9];
				11'd510:E2 <= line_E09[38];	11'd520:E2 <= line_E09[28];	11'd530:E2 <= line_E09[18];	11'd540:E2 <= line_E09[8];
				11'd511:E2 <= line_E09[37];	11'd521:E2 <= line_E09[27];	11'd531:E2 <= line_E09[17];	11'd541:E2 <= line_E09[7];
				11'd512:E2 <= line_E09[36];	11'd522:E2 <= line_E09[26];	11'd532:E2 <= line_E09[16];	11'd542:E2 <= line_E09[6];
				11'd513:E2 <= line_E09[35];	11'd523:E2 <= line_E09[25];	11'd533:E2 <= line_E09[15];	11'd543:E2 <= line_E09[5];
				11'd514:E2 <= line_E09[34];	11'd524:E2 <= line_E09[24];	11'd534:E2 <= line_E09[14];	11'd544:E2 <= line_E09[4];
				11'd515:E2 <= line_E09[33];	11'd525:E2 <= line_E09[23];	11'd535:E2 <= line_E09[13];	11'd545:E2 <= line_E09[3];
				11'd516:E2 <= line_E09[32];	11'd526:E2 <= line_E09[22];	11'd536:E2 <= line_E09[12];	11'd546:E2 <= line_E09[2];
				11'd517:E2 <= line_E09[31];	11'd527:E2 <= line_E09[21];	11'd537:E2 <= line_E09[11];	11'd547:E2 <= line_E09[1];
				11'd518:E2 <= line_E09[30];	11'd528:E2 <= line_E09[20];	11'd538:E2 <= line_E09[10];	11'd548:E2 <= line_E09[0];
				default:E2 <= 0;
			endcase
		11'd357:
			case (pixel_col)
				11'd509:E2 <= line_E10[39];	11'd519:E2 <= line_E10[29];	11'd529:E2 <= line_E10[19];	11'd539:E2 <= line_E10[9];
				11'd510:E2 <= line_E10[38];	11'd520:E2 <= line_E10[28];	11'd530:E2 <= line_E10[18];	11'd540:E2 <= line_E10[8];
				11'd511:E2 <= line_E10[37];	11'd521:E2 <= line_E10[27];	11'd531:E2 <= line_E10[17];	11'd541:E2 <= line_E10[7];
				11'd512:E2 <= line_E10[36];	11'd522:E2 <= line_E10[26];	11'd532:E2 <= line_E10[16];	11'd542:E2 <= line_E10[6];
				11'd513:E2 <= line_E10[35];	11'd523:E2 <= line_E10[25];	11'd533:E2 <= line_E10[15];	11'd543:E2 <= line_E10[5];
				11'd514:E2 <= line_E10[34];	11'd524:E2 <= line_E10[24];	11'd534:E2 <= line_E10[14];	11'd544:E2 <= line_E10[4];
				11'd515:E2 <= line_E10[33];	11'd525:E2 <= line_E10[23];	11'd535:E2 <= line_E10[13];	11'd545:E2 <= line_E10[3];
				11'd516:E2 <= line_E10[32];	11'd526:E2 <= line_E10[22];	11'd536:E2 <= line_E10[12];	11'd546:E2 <= line_E10[2];
				11'd517:E2 <= line_E10[31];	11'd527:E2 <= line_E10[21];	11'd537:E2 <= line_E10[11];	11'd547:E2 <= line_E10[1];
				11'd518:E2 <= line_E10[30];	11'd528:E2 <= line_E10[20];	11'd538:E2 <= line_E10[10];	11'd548:E2 <= line_E10[0];
				default:E2 <= 0;
			endcase
		11'd358:
			case (pixel_col)
				11'd509:E2 <= line_E11[39];	11'd519:E2 <= line_E11[29];	11'd529:E2 <= line_E11[19];	11'd539:E2 <= line_E11[9];
				11'd510:E2 <= line_E11[38];	11'd520:E2 <= line_E11[28];	11'd530:E2 <= line_E11[18];	11'd540:E2 <= line_E11[8];
				11'd511:E2 <= line_E11[37];	11'd521:E2 <= line_E11[27];	11'd531:E2 <= line_E11[17];	11'd541:E2 <= line_E11[7];
				11'd512:E2 <= line_E11[36];	11'd522:E2 <= line_E11[26];	11'd532:E2 <= line_E11[16];	11'd542:E2 <= line_E11[6];
				11'd513:E2 <= line_E11[35];	11'd523:E2 <= line_E11[25];	11'd533:E2 <= line_E11[15];	11'd543:E2 <= line_E11[5];
				11'd514:E2 <= line_E11[34];	11'd524:E2 <= line_E11[24];	11'd534:E2 <= line_E11[14];	11'd544:E2 <= line_E11[4];
				11'd515:E2 <= line_E11[33];	11'd525:E2 <= line_E11[23];	11'd535:E2 <= line_E11[13];	11'd545:E2 <= line_E11[3];
				11'd516:E2 <= line_E11[32];	11'd526:E2 <= line_E11[22];	11'd536:E2 <= line_E11[12];	11'd546:E2 <= line_E11[2];
				11'd517:E2 <= line_E11[31];	11'd527:E2 <= line_E11[21];	11'd537:E2 <= line_E11[11];	11'd547:E2 <= line_E11[1];
				11'd518:E2 <= line_E11[30];	11'd528:E2 <= line_E11[20];	11'd538:E2 <= line_E11[10];	11'd548:E2 <= line_E11[0];
				default:E2 <= 0;
			endcase
		11'd359:
			case (pixel_col)
				11'd509:E2 <= line_E12[39];	11'd519:E2 <= line_E12[29];	11'd529:E2 <= line_E12[19];	11'd539:E2 <= line_E12[9];
				11'd510:E2 <= line_E12[38];	11'd520:E2 <= line_E12[28];	11'd530:E2 <= line_E12[18];	11'd540:E2 <= line_E12[8];
				11'd511:E2 <= line_E12[37];	11'd521:E2 <= line_E12[27];	11'd531:E2 <= line_E12[17];	11'd541:E2 <= line_E12[7];
				11'd512:E2 <= line_E12[36];	11'd522:E2 <= line_E12[26];	11'd532:E2 <= line_E12[16];	11'd542:E2 <= line_E12[6];
				11'd513:E2 <= line_E12[35];	11'd523:E2 <= line_E12[25];	11'd533:E2 <= line_E12[15];	11'd543:E2 <= line_E12[5];
				11'd514:E2 <= line_E12[34];	11'd524:E2 <= line_E12[24];	11'd534:E2 <= line_E12[14];	11'd544:E2 <= line_E12[4];
				11'd515:E2 <= line_E12[33];	11'd525:E2 <= line_E12[23];	11'd535:E2 <= line_E12[13];	11'd545:E2 <= line_E12[3];
				11'd516:E2 <= line_E12[32];	11'd526:E2 <= line_E12[22];	11'd536:E2 <= line_E12[12];	11'd546:E2 <= line_E12[2];
				11'd517:E2 <= line_E12[31];	11'd527:E2 <= line_E12[21];	11'd537:E2 <= line_E12[11];	11'd547:E2 <= line_E12[1];
				11'd518:E2 <= line_E12[30];	11'd528:E2 <= line_E12[20];	11'd538:E2 <= line_E12[10];	11'd548:E2 <= line_E12[0];
				default:E2 <= 0;
			endcase
		11'd360:
			case (pixel_col)
				11'd509:E2 <= line_E13[39];	11'd519:E2 <= line_E13[29];	11'd529:E2 <= line_E13[19];	11'd539:E2 <= line_E13[9];
				11'd510:E2 <= line_E13[38];	11'd520:E2 <= line_E13[28];	11'd530:E2 <= line_E13[18];	11'd540:E2 <= line_E13[8];
				11'd511:E2 <= line_E13[37];	11'd521:E2 <= line_E13[27];	11'd531:E2 <= line_E13[17];	11'd541:E2 <= line_E13[7];
				11'd512:E2 <= line_E13[36];	11'd522:E2 <= line_E13[26];	11'd532:E2 <= line_E13[16];	11'd542:E2 <= line_E13[6];
				11'd513:E2 <= line_E13[35];	11'd523:E2 <= line_E13[25];	11'd533:E2 <= line_E13[15];	11'd543:E2 <= line_E13[5];
				11'd514:E2 <= line_E13[34];	11'd524:E2 <= line_E13[24];	11'd534:E2 <= line_E13[14];	11'd544:E2 <= line_E13[4];
				11'd515:E2 <= line_E13[33];	11'd525:E2 <= line_E13[23];	11'd535:E2 <= line_E13[13];	11'd545:E2 <= line_E13[3];
				11'd516:E2 <= line_E13[32];	11'd526:E2 <= line_E13[22];	11'd536:E2 <= line_E13[12];	11'd546:E2 <= line_E13[2];
				11'd517:E2 <= line_E13[31];	11'd527:E2 <= line_E13[21];	11'd537:E2 <= line_E13[11];	11'd547:E2 <= line_E13[1];
				11'd518:E2 <= line_E13[30];	11'd528:E2 <= line_E13[20];	11'd538:E2 <= line_E13[10];	11'd548:E2 <= line_E13[0];
				default:E2 <= 0;
			endcase
		11'd361:
			case (pixel_col)
				11'd509:E2 <= line_E14[39];	11'd519:E2 <= line_E14[29];	11'd529:E2 <= line_E14[19];	11'd539:E2 <= line_E14[9];
				11'd510:E2 <= line_E14[38];	11'd520:E2 <= line_E14[28];	11'd530:E2 <= line_E14[18];	11'd540:E2 <= line_E14[8];
				11'd511:E2 <= line_E14[37];	11'd521:E2 <= line_E14[27];	11'd531:E2 <= line_E14[17];	11'd541:E2 <= line_E14[7];
				11'd512:E2 <= line_E14[36];	11'd522:E2 <= line_E14[26];	11'd532:E2 <= line_E14[16];	11'd542:E2 <= line_E14[6];
				11'd513:E2 <= line_E14[35];	11'd523:E2 <= line_E14[25];	11'd533:E2 <= line_E14[15];	11'd543:E2 <= line_E14[5];
				11'd514:E2 <= line_E14[34];	11'd524:E2 <= line_E14[24];	11'd534:E2 <= line_E14[14];	11'd544:E2 <= line_E14[4];
				11'd515:E2 <= line_E14[33];	11'd525:E2 <= line_E14[23];	11'd535:E2 <= line_E14[13];	11'd545:E2 <= line_E14[3];
				11'd516:E2 <= line_E14[32];	11'd526:E2 <= line_E14[22];	11'd536:E2 <= line_E14[12];	11'd546:E2 <= line_E14[2];
				11'd517:E2 <= line_E14[31];	11'd527:E2 <= line_E14[21];	11'd537:E2 <= line_E14[11];	11'd547:E2 <= line_E14[1];
				11'd518:E2 <= line_E14[30];	11'd528:E2 <= line_E14[20];	11'd538:E2 <= line_E14[10];	11'd548:E2 <= line_E14[0];
				default:E2 <= 0;
			endcase
		11'd362:
			case (pixel_col)
				11'd509:E2 <= line_E15[39];	11'd519:E2 <= line_E15[29];	11'd529:E2 <= line_E15[19];	11'd539:E2 <= line_E15[9];
				11'd510:E2 <= line_E15[38];	11'd520:E2 <= line_E15[28];	11'd530:E2 <= line_E15[18];	11'd540:E2 <= line_E15[8];
				11'd511:E2 <= line_E15[37];	11'd521:E2 <= line_E15[27];	11'd531:E2 <= line_E15[17];	11'd541:E2 <= line_E15[7];
				11'd512:E2 <= line_E15[36];	11'd522:E2 <= line_E15[26];	11'd532:E2 <= line_E15[16];	11'd542:E2 <= line_E15[6];
				11'd513:E2 <= line_E15[35];	11'd523:E2 <= line_E15[25];	11'd533:E2 <= line_E15[15];	11'd543:E2 <= line_E15[5];
				11'd514:E2 <= line_E15[34];	11'd524:E2 <= line_E15[24];	11'd534:E2 <= line_E15[14];	11'd544:E2 <= line_E15[4];
				11'd515:E2 <= line_E15[33];	11'd525:E2 <= line_E15[23];	11'd535:E2 <= line_E15[13];	11'd545:E2 <= line_E15[3];
				11'd516:E2 <= line_E15[32];	11'd526:E2 <= line_E15[22];	11'd536:E2 <= line_E15[12];	11'd546:E2 <= line_E15[2];
				11'd517:E2 <= line_E15[31];	11'd527:E2 <= line_E15[21];	11'd537:E2 <= line_E15[11];	11'd547:E2 <= line_E15[1];
				11'd518:E2 <= line_E15[30];	11'd528:E2 <= line_E15[20];	11'd538:E2 <= line_E15[10];	11'd548:E2 <= line_E15[0];
				default:E2 <= 0;
			endcase
		default:E2 <= 0;
	endcase
end


always @(posedge clk) begin
	case (pixel_row)
		11'd348:
			case (pixel_col)
				11'd559:R <= line_R01[39];	11'd569:R <= line_R01[29];	11'd579:R <= line_R01[19];	11'd589:R <= line_R01[9];
				11'd560:R <= line_R01[38];	11'd570:R <= line_R01[28];	11'd580:R <= line_R01[18];	11'd590:R <= line_R01[8];
				11'd561:R <= line_R01[37];	11'd571:R <= line_R01[27];	11'd581:R <= line_R01[17];	11'd591:R <= line_R01[7];
				11'd562:R <= line_R01[36];	11'd572:R <= line_R01[26];	11'd582:R <= line_R01[16];	11'd592:R <= line_R01[6];
				11'd563:R <= line_R01[35];	11'd573:R <= line_R01[25];	11'd583:R <= line_R01[15];	11'd593:R <= line_R01[5];
				11'd564:R <= line_R01[34];	11'd574:R <= line_R01[24];	11'd584:R <= line_R01[14];	11'd594:R <= line_R01[4];
				11'd565:R <= line_R01[33];	11'd575:R <= line_R01[23];	11'd585:R <= line_R01[13];	11'd595:R <= line_R01[3];
				11'd566:R <= line_R01[32];	11'd576:R <= line_R01[22];	11'd586:R <= line_R01[12];	11'd596:R <= line_R01[2];
				11'd567:R <= line_R01[31];	11'd577:R <= line_R01[21];	11'd587:R <= line_R01[11];	11'd597:R <= line_R01[1];
				11'd568:R <= line_R01[30];	11'd578:R <= line_R01[20];	11'd588:R <= line_R01[10];	11'd598:R <= line_R01[0];
				default:R <= 0;
			endcase
		11'd349:
			case (pixel_col)
				11'd559:R <= line_R02[39];	11'd569:R <= line_R02[29];	11'd579:R <= line_R02[19];	11'd589:R <= line_R02[9];
				11'd560:R <= line_R02[38];	11'd570:R <= line_R02[28];	11'd580:R <= line_R02[18];	11'd590:R <= line_R02[8];
				11'd561:R <= line_R02[37];	11'd571:R <= line_R02[27];	11'd581:R <= line_R02[17];	11'd591:R <= line_R02[7];
				11'd562:R <= line_R02[36];	11'd572:R <= line_R02[26];	11'd582:R <= line_R02[16];	11'd592:R <= line_R02[6];
				11'd563:R <= line_R02[35];	11'd573:R <= line_R02[25];	11'd583:R <= line_R02[15];	11'd593:R <= line_R02[5];
				11'd564:R <= line_R02[34];	11'd574:R <= line_R02[24];	11'd584:R <= line_R02[14];	11'd594:R <= line_R02[4];
				11'd565:R <= line_R02[33];	11'd575:R <= line_R02[23];	11'd585:R <= line_R02[13];	11'd595:R <= line_R02[3];
				11'd566:R <= line_R02[32];	11'd576:R <= line_R02[22];	11'd586:R <= line_R02[12];	11'd596:R <= line_R02[2];
				11'd567:R <= line_R02[31];	11'd577:R <= line_R02[21];	11'd587:R <= line_R02[11];	11'd597:R <= line_R02[1];
				11'd568:R <= line_R02[30];	11'd578:R <= line_R02[20];	11'd588:R <= line_R02[10];	11'd598:R <= line_R02[0];
				default:R <= 0;
			endcase
		11'd350:
			case (pixel_col)
				11'd559:R <= line_R03[39];	11'd569:R <= line_R03[29];	11'd579:R <= line_R03[19];	11'd589:R <= line_R03[9];
				11'd560:R <= line_R03[38];	11'd570:R <= line_R03[28];	11'd580:R <= line_R03[18];	11'd590:R <= line_R03[8];
				11'd561:R <= line_R03[37];	11'd571:R <= line_R03[27];	11'd581:R <= line_R03[17];	11'd591:R <= line_R03[7];
				11'd562:R <= line_R03[36];	11'd572:R <= line_R03[26];	11'd582:R <= line_R03[16];	11'd592:R <= line_R03[6];
				11'd563:R <= line_R03[35];	11'd573:R <= line_R03[25];	11'd583:R <= line_R03[15];	11'd593:R <= line_R03[5];
				11'd564:R <= line_R03[34];	11'd574:R <= line_R03[24];	11'd584:R <= line_R03[14];	11'd594:R <= line_R03[4];
				11'd565:R <= line_R03[33];	11'd575:R <= line_R03[23];	11'd585:R <= line_R03[13];	11'd595:R <= line_R03[3];
				11'd566:R <= line_R03[32];	11'd576:R <= line_R03[22];	11'd586:R <= line_R03[12];	11'd596:R <= line_R03[2];
				11'd567:R <= line_R03[31];	11'd577:R <= line_R03[21];	11'd587:R <= line_R03[11];	11'd597:R <= line_R03[1];
				11'd568:R <= line_R03[30];	11'd578:R <= line_R03[20];	11'd588:R <= line_R03[10];	11'd598:R <= line_R03[0];
				default:R <= 0;
			endcase
		11'd351:
			case (pixel_col)
				11'd559:R <= line_R04[39];	11'd569:R <= line_R04[29];	11'd579:R <= line_R04[19];	11'd589:R <= line_R04[9];
				11'd560:R <= line_R04[38];	11'd570:R <= line_R04[28];	11'd580:R <= line_R04[18];	11'd590:R <= line_R04[8];
				11'd561:R <= line_R04[37];	11'd571:R <= line_R04[27];	11'd581:R <= line_R04[17];	11'd591:R <= line_R04[7];
				11'd562:R <= line_R04[36];	11'd572:R <= line_R04[26];	11'd582:R <= line_R04[16];	11'd592:R <= line_R04[6];
				11'd563:R <= line_R04[35];	11'd573:R <= line_R04[25];	11'd583:R <= line_R04[15];	11'd593:R <= line_R04[5];
				11'd564:R <= line_R04[34];	11'd574:R <= line_R04[24];	11'd584:R <= line_R04[14];	11'd594:R <= line_R04[4];
				11'd565:R <= line_R04[33];	11'd575:R <= line_R04[23];	11'd585:R <= line_R04[13];	11'd595:R <= line_R04[3];
				11'd566:R <= line_R04[32];	11'd576:R <= line_R04[22];	11'd586:R <= line_R04[12];	11'd596:R <= line_R04[2];
				11'd567:R <= line_R04[31];	11'd577:R <= line_R04[21];	11'd587:R <= line_R04[11];	11'd597:R <= line_R04[1];
				11'd568:R <= line_R04[30];	11'd578:R <= line_R04[20];	11'd588:R <= line_R04[10];	11'd598:R <= line_R04[0];
				default:R <= 0;
			endcase
		11'd352:
			case (pixel_col)
				11'd559:R <= line_R05[39];	11'd569:R <= line_R05[29];	11'd579:R <= line_R05[19];	11'd589:R <= line_R05[9];
				11'd560:R <= line_R05[38];	11'd570:R <= line_R05[28];	11'd580:R <= line_R05[18];	11'd590:R <= line_R05[8];
				11'd561:R <= line_R05[37];	11'd571:R <= line_R05[27];	11'd581:R <= line_R05[17];	11'd591:R <= line_R05[7];
				11'd562:R <= line_R05[36];	11'd572:R <= line_R05[26];	11'd582:R <= line_R05[16];	11'd592:R <= line_R05[6];
				11'd563:R <= line_R05[35];	11'd573:R <= line_R05[25];	11'd583:R <= line_R05[15];	11'd593:R <= line_R05[5];
				11'd564:R <= line_R05[34];	11'd574:R <= line_R05[24];	11'd584:R <= line_R05[14];	11'd594:R <= line_R05[4];
				11'd565:R <= line_R05[33];	11'd575:R <= line_R05[23];	11'd585:R <= line_R05[13];	11'd595:R <= line_R05[3];
				11'd566:R <= line_R05[32];	11'd576:R <= line_R05[22];	11'd586:R <= line_R05[12];	11'd596:R <= line_R05[2];
				11'd567:R <= line_R05[31];	11'd577:R <= line_R05[21];	11'd587:R <= line_R05[11];	11'd597:R <= line_R05[1];
				11'd568:R <= line_R05[30];	11'd578:R <= line_R05[20];	11'd588:R <= line_R05[10];	11'd598:R <= line_R05[0];
				default:R <= 0;
			endcase
		11'd353:
			case (pixel_col)
				11'd559:R <= line_R06[39];	11'd569:R <= line_R06[29];	11'd579:R <= line_R06[19];	11'd589:R <= line_R06[9];
				11'd560:R <= line_R06[38];	11'd570:R <= line_R06[28];	11'd580:R <= line_R06[18];	11'd590:R <= line_R06[8];
				11'd561:R <= line_R06[37];	11'd571:R <= line_R06[27];	11'd581:R <= line_R06[17];	11'd591:R <= line_R06[7];
				11'd562:R <= line_R06[36];	11'd572:R <= line_R06[26];	11'd582:R <= line_R06[16];	11'd592:R <= line_R06[6];
				11'd563:R <= line_R06[35];	11'd573:R <= line_R06[25];	11'd583:R <= line_R06[15];	11'd593:R <= line_R06[5];
				11'd564:R <= line_R06[34];	11'd574:R <= line_R06[24];	11'd584:R <= line_R06[14];	11'd594:R <= line_R06[4];
				11'd565:R <= line_R06[33];	11'd575:R <= line_R06[23];	11'd585:R <= line_R06[13];	11'd595:R <= line_R06[3];
				11'd566:R <= line_R06[32];	11'd576:R <= line_R06[22];	11'd586:R <= line_R06[12];	11'd596:R <= line_R06[2];
				11'd567:R <= line_R06[31];	11'd577:R <= line_R06[21];	11'd587:R <= line_R06[11];	11'd597:R <= line_R06[1];
				11'd568:R <= line_R06[30];	11'd578:R <= line_R06[20];	11'd588:R <= line_R06[10];	11'd598:R <= line_R06[0];
				default:R <= 0;
			endcase
		11'd354:
			case (pixel_col)
				11'd559:R <= line_R07[39];	11'd569:R <= line_R07[29];	11'd579:R <= line_R07[19];	11'd589:R <= line_R07[9];
				11'd560:R <= line_R07[38];	11'd570:R <= line_R07[28];	11'd580:R <= line_R07[18];	11'd590:R <= line_R07[8];
				11'd561:R <= line_R07[37];	11'd571:R <= line_R07[27];	11'd581:R <= line_R07[17];	11'd591:R <= line_R07[7];
				11'd562:R <= line_R07[36];	11'd572:R <= line_R07[26];	11'd582:R <= line_R07[16];	11'd592:R <= line_R07[6];
				11'd563:R <= line_R07[35];	11'd573:R <= line_R07[25];	11'd583:R <= line_R07[15];	11'd593:R <= line_R07[5];
				11'd564:R <= line_R07[34];	11'd574:R <= line_R07[24];	11'd584:R <= line_R07[14];	11'd594:R <= line_R07[4];
				11'd565:R <= line_R07[33];	11'd575:R <= line_R07[23];	11'd585:R <= line_R07[13];	11'd595:R <= line_R07[3];
				11'd566:R <= line_R07[32];	11'd576:R <= line_R07[22];	11'd586:R <= line_R07[12];	11'd596:R <= line_R07[2];
				11'd567:R <= line_R07[31];	11'd577:R <= line_R07[21];	11'd587:R <= line_R07[11];	11'd597:R <= line_R07[1];
				11'd568:R <= line_R07[30];	11'd578:R <= line_R07[20];	11'd588:R <= line_R07[10];	11'd598:R <= line_R07[0];
				default:R <= 0;
			endcase
		11'd355:
			case (pixel_col)
				11'd559:R <= line_R08[39];	11'd569:R <= line_R08[29];	11'd579:R <= line_R08[19];	11'd589:R <= line_R08[9];
				11'd560:R <= line_R08[38];	11'd570:R <= line_R08[28];	11'd580:R <= line_R08[18];	11'd590:R <= line_R08[8];
				11'd561:R <= line_R08[37];	11'd571:R <= line_R08[27];	11'd581:R <= line_R08[17];	11'd591:R <= line_R08[7];
				11'd562:R <= line_R08[36];	11'd572:R <= line_R08[26];	11'd582:R <= line_R08[16];	11'd592:R <= line_R08[6];
				11'd563:R <= line_R08[35];	11'd573:R <= line_R08[25];	11'd583:R <= line_R08[15];	11'd593:R <= line_R08[5];
				11'd564:R <= line_R08[34];	11'd574:R <= line_R08[24];	11'd584:R <= line_R08[14];	11'd594:R <= line_R08[4];
				11'd565:R <= line_R08[33];	11'd575:R <= line_R08[23];	11'd585:R <= line_R08[13];	11'd595:R <= line_R08[3];
				11'd566:R <= line_R08[32];	11'd576:R <= line_R08[22];	11'd586:R <= line_R08[12];	11'd596:R <= line_R08[2];
				11'd567:R <= line_R08[31];	11'd577:R <= line_R08[21];	11'd587:R <= line_R08[11];	11'd597:R <= line_R08[1];
				11'd568:R <= line_R08[30];	11'd578:R <= line_R08[20];	11'd588:R <= line_R08[10];	11'd598:R <= line_R08[0];
				default:R <= 0;
			endcase
		11'd356:
			case (pixel_col)
				11'd559:R <= line_R09[39];	11'd569:R <= line_R09[29];	11'd579:R <= line_R09[19];	11'd589:R <= line_R09[9];
				11'd560:R <= line_R09[38];	11'd570:R <= line_R09[28];	11'd580:R <= line_R09[18];	11'd590:R <= line_R09[8];
				11'd561:R <= line_R09[37];	11'd571:R <= line_R09[27];	11'd581:R <= line_R09[17];	11'd591:R <= line_R09[7];
				11'd562:R <= line_R09[36];	11'd572:R <= line_R09[26];	11'd582:R <= line_R09[16];	11'd592:R <= line_R09[6];
				11'd563:R <= line_R09[35];	11'd573:R <= line_R09[25];	11'd583:R <= line_R09[15];	11'd593:R <= line_R09[5];
				11'd564:R <= line_R09[34];	11'd574:R <= line_R09[24];	11'd584:R <= line_R09[14];	11'd594:R <= line_R09[4];
				11'd565:R <= line_R09[33];	11'd575:R <= line_R09[23];	11'd585:R <= line_R09[13];	11'd595:R <= line_R09[3];
				11'd566:R <= line_R09[32];	11'd576:R <= line_R09[22];	11'd586:R <= line_R09[12];	11'd596:R <= line_R09[2];
				11'd567:R <= line_R09[31];	11'd577:R <= line_R09[21];	11'd587:R <= line_R09[11];	11'd597:R <= line_R09[1];
				11'd568:R <= line_R09[30];	11'd578:R <= line_R09[20];	11'd588:R <= line_R09[10];	11'd598:R <= line_R09[0];
				default:R <= 0;
			endcase
		11'd357:
			case (pixel_col)
				11'd559:R <= line_R10[39];	11'd569:R <= line_R10[29];	11'd579:R <= line_R10[19];	11'd589:R <= line_R10[9];
				11'd560:R <= line_R10[38];	11'd570:R <= line_R10[28];	11'd580:R <= line_R10[18];	11'd590:R <= line_R10[8];
				11'd561:R <= line_R10[37];	11'd571:R <= line_R10[27];	11'd581:R <= line_R10[17];	11'd591:R <= line_R10[7];
				11'd562:R <= line_R10[36];	11'd572:R <= line_R10[26];	11'd582:R <= line_R10[16];	11'd592:R <= line_R10[6];
				11'd563:R <= line_R10[35];	11'd573:R <= line_R10[25];	11'd583:R <= line_R10[15];	11'd593:R <= line_R10[5];
				11'd564:R <= line_R10[34];	11'd574:R <= line_R10[24];	11'd584:R <= line_R10[14];	11'd594:R <= line_R10[4];
				11'd565:R <= line_R10[33];	11'd575:R <= line_R10[23];	11'd585:R <= line_R10[13];	11'd595:R <= line_R10[3];
				11'd566:R <= line_R10[32];	11'd576:R <= line_R10[22];	11'd586:R <= line_R10[12];	11'd596:R <= line_R10[2];
				11'd567:R <= line_R10[31];	11'd577:R <= line_R10[21];	11'd587:R <= line_R10[11];	11'd597:R <= line_R10[1];
				11'd568:R <= line_R10[30];	11'd578:R <= line_R10[20];	11'd588:R <= line_R10[10];	11'd598:R <= line_R10[0];
				default:R <= 0;
			endcase
		11'd358:
			case (pixel_col)
				11'd559:R <= line_R11[39];	11'd569:R <= line_R11[29];	11'd579:R <= line_R11[19];	11'd589:R <= line_R11[9];
				11'd560:R <= line_R11[38];	11'd570:R <= line_R11[28];	11'd580:R <= line_R11[18];	11'd590:R <= line_R11[8];
				11'd561:R <= line_R11[37];	11'd571:R <= line_R11[27];	11'd581:R <= line_R11[17];	11'd591:R <= line_R11[7];
				11'd562:R <= line_R11[36];	11'd572:R <= line_R11[26];	11'd582:R <= line_R11[16];	11'd592:R <= line_R11[6];
				11'd563:R <= line_R11[35];	11'd573:R <= line_R11[25];	11'd583:R <= line_R11[15];	11'd593:R <= line_R11[5];
				11'd564:R <= line_R11[34];	11'd574:R <= line_R11[24];	11'd584:R <= line_R11[14];	11'd594:R <= line_R11[4];
				11'd565:R <= line_R11[33];	11'd575:R <= line_R11[23];	11'd585:R <= line_R11[13];	11'd595:R <= line_R11[3];
				11'd566:R <= line_R11[32];	11'd576:R <= line_R11[22];	11'd586:R <= line_R11[12];	11'd596:R <= line_R11[2];
				11'd567:R <= line_R11[31];	11'd577:R <= line_R11[21];	11'd587:R <= line_R11[11];	11'd597:R <= line_R11[1];
				11'd568:R <= line_R11[30];	11'd578:R <= line_R11[20];	11'd588:R <= line_R11[10];	11'd598:R <= line_R11[0];
				default:R <= 0;
			endcase
		11'd359:
			case (pixel_col)
				11'd559:R <= line_R12[39];	11'd569:R <= line_R12[29];	11'd579:R <= line_R12[19];	11'd589:R <= line_R12[9];
				11'd560:R <= line_R12[38];	11'd570:R <= line_R12[28];	11'd580:R <= line_R12[18];	11'd590:R <= line_R12[8];
				11'd561:R <= line_R12[37];	11'd571:R <= line_R12[27];	11'd581:R <= line_R12[17];	11'd591:R <= line_R12[7];
				11'd562:R <= line_R12[36];	11'd572:R <= line_R12[26];	11'd582:R <= line_R12[16];	11'd592:R <= line_R12[6];
				11'd563:R <= line_R12[35];	11'd573:R <= line_R12[25];	11'd583:R <= line_R12[15];	11'd593:R <= line_R12[5];
				11'd564:R <= line_R12[34];	11'd574:R <= line_R12[24];	11'd584:R <= line_R12[14];	11'd594:R <= line_R12[4];
				11'd565:R <= line_R12[33];	11'd575:R <= line_R12[23];	11'd585:R <= line_R12[13];	11'd595:R <= line_R12[3];
				11'd566:R <= line_R12[32];	11'd576:R <= line_R12[22];	11'd586:R <= line_R12[12];	11'd596:R <= line_R12[2];
				11'd567:R <= line_R12[31];	11'd577:R <= line_R12[21];	11'd587:R <= line_R12[11];	11'd597:R <= line_R12[1];
				11'd568:R <= line_R12[30];	11'd578:R <= line_R12[20];	11'd588:R <= line_R12[10];	11'd598:R <= line_R12[0];
				default:R <= 0;
			endcase
		11'd360:
			case (pixel_col)
				11'd559:R <= line_R13[39];	11'd569:R <= line_R13[29];	11'd579:R <= line_R13[19];	11'd589:R <= line_R13[9];
				11'd560:R <= line_R13[38];	11'd570:R <= line_R13[28];	11'd580:R <= line_R13[18];	11'd590:R <= line_R13[8];
				11'd561:R <= line_R13[37];	11'd571:R <= line_R13[27];	11'd581:R <= line_R13[17];	11'd591:R <= line_R13[7];
				11'd562:R <= line_R13[36];	11'd572:R <= line_R13[26];	11'd582:R <= line_R13[16];	11'd592:R <= line_R13[6];
				11'd563:R <= line_R13[35];	11'd573:R <= line_R13[25];	11'd583:R <= line_R13[15];	11'd593:R <= line_R13[5];
				11'd564:R <= line_R13[34];	11'd574:R <= line_R13[24];	11'd584:R <= line_R13[14];	11'd594:R <= line_R13[4];
				11'd565:R <= line_R13[33];	11'd575:R <= line_R13[23];	11'd585:R <= line_R13[13];	11'd595:R <= line_R13[3];
				11'd566:R <= line_R13[32];	11'd576:R <= line_R13[22];	11'd586:R <= line_R13[12];	11'd596:R <= line_R13[2];
				11'd567:R <= line_R13[31];	11'd577:R <= line_R13[21];	11'd587:R <= line_R13[11];	11'd597:R <= line_R13[1];
				11'd568:R <= line_R13[30];	11'd578:R <= line_R13[20];	11'd588:R <= line_R13[10];	11'd598:R <= line_R13[0];
				default:R <= 0;
			endcase
		11'd361:
			case (pixel_col)
				11'd559:R <= line_R14[39];	11'd569:R <= line_R14[29];	11'd579:R <= line_R14[19];	11'd589:R <= line_R14[9];
				11'd560:R <= line_R14[38];	11'd570:R <= line_R14[28];	11'd580:R <= line_R14[18];	11'd590:R <= line_R14[8];
				11'd561:R <= line_R14[37];	11'd571:R <= line_R14[27];	11'd581:R <= line_R14[17];	11'd591:R <= line_R14[7];
				11'd562:R <= line_R14[36];	11'd572:R <= line_R14[26];	11'd582:R <= line_R14[16];	11'd592:R <= line_R14[6];
				11'd563:R <= line_R14[35];	11'd573:R <= line_R14[25];	11'd583:R <= line_R14[15];	11'd593:R <= line_R14[5];
				11'd564:R <= line_R14[34];	11'd574:R <= line_R14[24];	11'd584:R <= line_R14[14];	11'd594:R <= line_R14[4];
				11'd565:R <= line_R14[33];	11'd575:R <= line_R14[23];	11'd585:R <= line_R14[13];	11'd595:R <= line_R14[3];
				11'd566:R <= line_R14[32];	11'd576:R <= line_R14[22];	11'd586:R <= line_R14[12];	11'd596:R <= line_R14[2];
				11'd567:R <= line_R14[31];	11'd577:R <= line_R14[21];	11'd587:R <= line_R14[11];	11'd597:R <= line_R14[1];
				11'd568:R <= line_R14[30];	11'd578:R <= line_R14[20];	11'd588:R <= line_R14[10];	11'd598:R <= line_R14[0];
				default:R <= 0;
			endcase
		11'd362:
			case (pixel_col)
				11'd559:R <= line_R15[39];	11'd569:R <= line_R15[29];	11'd579:R <= line_R15[19];	11'd589:R <= line_R15[9];
				11'd560:R <= line_R15[38];	11'd570:R <= line_R15[28];	11'd580:R <= line_R15[18];	11'd590:R <= line_R15[8];
				11'd561:R <= line_R15[37];	11'd571:R <= line_R15[27];	11'd581:R <= line_R15[17];	11'd591:R <= line_R15[7];
				11'd562:R <= line_R15[36];	11'd572:R <= line_R15[26];	11'd582:R <= line_R15[16];	11'd592:R <= line_R15[6];
				11'd563:R <= line_R15[35];	11'd573:R <= line_R15[25];	11'd583:R <= line_R15[15];	11'd593:R <= line_R15[5];
				11'd564:R <= line_R15[34];	11'd574:R <= line_R15[24];	11'd584:R <= line_R15[14];	11'd594:R <= line_R15[4];
				11'd565:R <= line_R15[33];	11'd575:R <= line_R15[23];	11'd585:R <= line_R15[13];	11'd595:R <= line_R15[3];
				11'd566:R <= line_R15[32];	11'd576:R <= line_R15[22];	11'd586:R <= line_R15[12];	11'd596:R <= line_R15[2];
				11'd567:R <= line_R15[31];	11'd577:R <= line_R15[21];	11'd587:R <= line_R15[11];	11'd597:R <= line_R15[1];
				11'd568:R <= line_R15[30];	11'd578:R <= line_R15[20];	11'd588:R <= line_R15[10];	11'd598:R <= line_R15[0];
				default:R <= 0;
			endcase
		default:R <= 0;
	endcase
end

endmodule 